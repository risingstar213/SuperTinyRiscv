module Core(
  input         clock,
  input         reset,
  output [31:0] io_imem_addr,
  input  [31:0] io_imem_inst,
  output [31:0] io_dmem_addr,
  input  [31:0] io_dmem_rdata,
  output        io_dmem_wen,
  output [31:0] io_dmem_wdata,
  output [2:0]  io_dmem_rwtype,
  output [31:0] io_data
);
  reg [31:0] regfile [0:31]; // @[Core.scala 17:22]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_8_data; // @[Core.scala 17:22]
  wire [4:0] regfile__T_8_addr; // @[Core.scala 17:22]
  wire [31:0] regfile__T_11_data; // @[Core.scala 17:22]
  wire [4:0] regfile__T_11_addr; // @[Core.scala 17:22]
  wire [31:0] regfile__T_18_data; // @[Core.scala 17:22]
  wire [4:0] regfile__T_18_addr; // @[Core.scala 17:22]
  wire [31:0] regfile__T_21_data; // @[Core.scala 17:22]
  wire [4:0] regfile__T_21_addr; // @[Core.scala 17:22]
  wire [31:0] regfile__T_568_data; // @[Core.scala 17:22]
  wire [4:0] regfile__T_568_addr; // @[Core.scala 17:22]
  wire  regfile__T_568_mask; // @[Core.scala 17:22]
  wire  regfile__T_568_en; // @[Core.scala 17:22]
  reg [31:0] pc_reg; // @[Core.scala 21:25]
  reg [31:0] _RAND_1;
  wire [31:0] pc_plus4; // @[Core.scala 25:27]
  wire [31:0] _T_1; // @[Core.scala 33:15]
  wire  _T_2; // @[Core.scala 33:15]
  wire [31:0] _T_3; // @[Core.scala 33:31]
  wire  _T_4; // @[Core.scala 33:31]
  wire  _T_5; // @[Core.scala 33:23]
  wire  _T_58; // @[Lookup.scala 31:38]
  wire  _T_60; // @[Lookup.scala 31:38]
  wire  _T_62; // @[Lookup.scala 31:38]
  wire  _T_64; // @[Lookup.scala 31:38]
  wire  _T_66; // @[Lookup.scala 31:38]
  wire  _T_68; // @[Lookup.scala 31:38]
  wire  _T_70; // @[Lookup.scala 31:38]
  wire  _T_72; // @[Lookup.scala 31:38]
  wire [31:0] _T_73; // @[Lookup.scala 31:38]
  wire  _T_74; // @[Lookup.scala 31:38]
  wire  _T_76; // @[Lookup.scala 31:38]
  wire  _T_78; // @[Lookup.scala 31:38]
  wire  _T_80; // @[Lookup.scala 31:38]
  wire  _T_82; // @[Lookup.scala 31:38]
  wire  _T_84; // @[Lookup.scala 31:38]
  wire  _T_86; // @[Lookup.scala 31:38]
  wire  _T_88; // @[Lookup.scala 31:38]
  wire  _T_90; // @[Lookup.scala 31:38]
  wire  _T_92; // @[Lookup.scala 31:38]
  wire  _T_94; // @[Lookup.scala 31:38]
  wire  _T_96; // @[Lookup.scala 31:38]
  wire  _T_98; // @[Lookup.scala 31:38]
  wire  _T_100; // @[Lookup.scala 31:38]
  wire  _T_102; // @[Lookup.scala 31:38]
  wire  _T_104; // @[Lookup.scala 31:38]
  wire  _T_106; // @[Lookup.scala 31:38]
  wire  _T_108; // @[Lookup.scala 31:38]
  wire  _T_110; // @[Lookup.scala 31:38]
  wire  _T_112; // @[Lookup.scala 31:38]
  wire  _T_114; // @[Lookup.scala 31:38]
  wire  _T_116; // @[Lookup.scala 31:38]
  wire  _T_118; // @[Lookup.scala 31:38]
  wire  _T_120; // @[Lookup.scala 31:38]
  wire  _T_122; // @[Lookup.scala 31:38]
  wire  _T_124; // @[Lookup.scala 31:38]
  wire  _T_126; // @[Lookup.scala 31:38]
  wire  _T_128; // @[Lookup.scala 31:38]
  wire  _T_130; // @[Lookup.scala 31:38]
  wire  _T_132; // @[Lookup.scala 31:38]
  wire  _T_134; // @[Lookup.scala 31:38]
  wire  _T_140; // @[Lookup.scala 31:38]
  wire  _T_142; // @[Lookup.scala 31:38]
  wire  _T_144; // @[Lookup.scala 31:38]
  wire [4:0] _T_145; // @[Lookup.scala 33:37]
  wire [4:0] _T_146; // @[Lookup.scala 33:37]
  wire [4:0] _T_147; // @[Lookup.scala 33:37]
  wire [4:0] _T_148; // @[Lookup.scala 33:37]
  wire [4:0] _T_149; // @[Lookup.scala 33:37]
  wire [4:0] _T_150; // @[Lookup.scala 33:37]
  wire [4:0] _T_151; // @[Lookup.scala 33:37]
  wire [4:0] _T_152; // @[Lookup.scala 33:37]
  wire [4:0] _T_153; // @[Lookup.scala 33:37]
  wire [4:0] _T_154; // @[Lookup.scala 33:37]
  wire [4:0] _T_155; // @[Lookup.scala 33:37]
  wire [4:0] _T_156; // @[Lookup.scala 33:37]
  wire [4:0] _T_157; // @[Lookup.scala 33:37]
  wire [4:0] _T_158; // @[Lookup.scala 33:37]
  wire [4:0] _T_159; // @[Lookup.scala 33:37]
  wire [4:0] _T_160; // @[Lookup.scala 33:37]
  wire [4:0] _T_161; // @[Lookup.scala 33:37]
  wire [4:0] _T_162; // @[Lookup.scala 33:37]
  wire [4:0] _T_163; // @[Lookup.scala 33:37]
  wire [4:0] _T_164; // @[Lookup.scala 33:37]
  wire [4:0] _T_165; // @[Lookup.scala 33:37]
  wire [4:0] _T_166; // @[Lookup.scala 33:37]
  wire [4:0] _T_167; // @[Lookup.scala 33:37]
  wire [4:0] _T_168; // @[Lookup.scala 33:37]
  wire [4:0] _T_169; // @[Lookup.scala 33:37]
  wire [4:0] _T_170; // @[Lookup.scala 33:37]
  wire [4:0] _T_171; // @[Lookup.scala 33:37]
  wire [4:0] _T_172; // @[Lookup.scala 33:37]
  wire [4:0] _T_173; // @[Lookup.scala 33:37]
  wire [4:0] _T_174; // @[Lookup.scala 33:37]
  wire [4:0] _T_175; // @[Lookup.scala 33:37]
  wire [4:0] _T_176; // @[Lookup.scala 33:37]
  wire [4:0] _T_177; // @[Lookup.scala 33:37]
  wire [4:0] _T_178; // @[Lookup.scala 33:37]
  wire [4:0] _T_179; // @[Lookup.scala 33:37]
  wire [4:0] _T_180; // @[Lookup.scala 33:37]
  wire [4:0] _T_181; // @[Lookup.scala 33:37]
  wire [4:0] _T_182; // @[Lookup.scala 33:37]
  wire [4:0] _T_183; // @[Lookup.scala 33:37]
  wire [4:0] _T_184; // @[Lookup.scala 33:37]
  wire [4:0] _T_185; // @[Lookup.scala 33:37]
  wire [4:0] _T_186; // @[Lookup.scala 33:37]
  wire [4:0] _T_187; // @[Lookup.scala 33:37]
  wire [4:0] csignals_0; // @[Lookup.scala 33:37]
  wire  _T_557; // @[Core.scala 163:27]
  wire [2:0] _T_232; // @[Lookup.scala 33:37]
  wire [2:0] _T_233; // @[Lookup.scala 33:37]
  wire [2:0] _T_234; // @[Lookup.scala 33:37]
  wire [2:0] _T_235; // @[Lookup.scala 33:37]
  wire [2:0] _T_236; // @[Lookup.scala 33:37]
  wire [2:0] _T_237; // @[Lookup.scala 33:37]
  wire [2:0] _T_238; // @[Lookup.scala 33:37]
  wire [2:0] _T_239; // @[Lookup.scala 33:37]
  wire [2:0] _T_240; // @[Lookup.scala 33:37]
  wire [2:0] _T_241; // @[Lookup.scala 33:37]
  wire [2:0] _T_242; // @[Lookup.scala 33:37]
  wire [2:0] _T_243; // @[Lookup.scala 33:37]
  wire [2:0] _T_244; // @[Lookup.scala 33:37]
  wire [2:0] _T_245; // @[Lookup.scala 33:37]
  wire [2:0] _T_246; // @[Lookup.scala 33:37]
  wire [2:0] _T_247; // @[Lookup.scala 33:37]
  wire [2:0] _T_248; // @[Lookup.scala 33:37]
  wire [2:0] _T_249; // @[Lookup.scala 33:37]
  wire [2:0] _T_250; // @[Lookup.scala 33:37]
  wire [2:0] _T_251; // @[Lookup.scala 33:37]
  wire [2:0] _T_252; // @[Lookup.scala 33:37]
  wire [2:0] _T_253; // @[Lookup.scala 33:37]
  wire [2:0] _T_254; // @[Lookup.scala 33:37]
  wire [2:0] _T_255; // @[Lookup.scala 33:37]
  wire [2:0] _T_256; // @[Lookup.scala 33:37]
  wire [2:0] _T_257; // @[Lookup.scala 33:37]
  wire [2:0] _T_258; // @[Lookup.scala 33:37]
  wire [2:0] _T_259; // @[Lookup.scala 33:37]
  wire [2:0] _T_260; // @[Lookup.scala 33:37]
  wire [2:0] _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_262; // @[Lookup.scala 33:37]
  wire [2:0] _T_263; // @[Lookup.scala 33:37]
  wire [2:0] _T_264; // @[Lookup.scala 33:37]
  wire [2:0] _T_265; // @[Lookup.scala 33:37]
  wire [2:0] _T_266; // @[Lookup.scala 33:37]
  wire [2:0] _T_267; // @[Lookup.scala 33:37]
  wire [2:0] _T_268; // @[Lookup.scala 33:37]
  wire [2:0] _T_269; // @[Lookup.scala 33:37]
  wire [2:0] _T_270; // @[Lookup.scala 33:37]
  wire [2:0] _T_271; // @[Lookup.scala 33:37]
  wire [2:0] _T_272; // @[Lookup.scala 33:37]
  wire [2:0] _T_273; // @[Lookup.scala 33:37]
  wire [2:0] csignals_2; // @[Lookup.scala 33:37]
  wire  _T_449; // @[Core.scala 122:18]
  wire  _T_24; // @[Core.scala 50:15]
  wire [4:0] rs2_addr; // @[Core.scala 41:24]
  wire  _T_25; // @[Core.scala 50:37]
  wire  _T_26; // @[Core.scala 50:25]
  wire [31:0] _T_27; // @[Mux.scala 87:16]
  wire [31:0] rs2_data; // @[Mux.scala 87:16]
  wire  _T_450; // @[Core.scala 123:18]
  wire [11:0] imm_i; // @[Core.scala 53:21]
  wire  _T_28; // @[Core.scala 54:40]
  wire [19:0] _T_30; // @[Bitwise.scala 71:12]
  wire [31:0] imm_i_sext; // @[Cat.scala 29:58]
  wire  _T_451; // @[Core.scala 124:18]
  wire [6:0] _T_31; // @[Core.scala 55:25]
  wire [4:0] _T_32; // @[Core.scala 55:39]
  wire [11:0] imm_s; // @[Cat.scala 29:58]
  wire  _T_33; // @[Core.scala 56:40]
  wire [19:0] _T_35; // @[Bitwise.scala 71:12]
  wire [31:0] imm_s_sext; // @[Cat.scala 29:58]
  wire  _T_452; // @[Core.scala 125:18]
  wire  _T_46; // @[Core.scala 59:25]
  wire [7:0] _T_47; // @[Core.scala 59:35]
  wire  _T_48; // @[Core.scala 59:49]
  wire [9:0] _T_49; // @[Core.scala 59:59]
  wire [19:0] imm_j; // @[Cat.scala 29:58]
  wire  _T_52; // @[Core.scala 60:40]
  wire [10:0] _T_54; // @[Bitwise.scala 71:12]
  wire [31:0] imm_j_sext; // @[Cat.scala 29:58]
  wire  _T_453; // @[Core.scala 126:18]
  wire [19:0] imm_u; // @[Core.scala 61:21]
  wire [31:0] imm_u_shifted; // @[Cat.scala 29:58]
  wire [31:0] _T_454; // @[Mux.scala 87:16]
  wire [31:0] _T_455; // @[Mux.scala 87:16]
  wire [31:0] _T_456; // @[Mux.scala 87:16]
  wire [31:0] _T_457; // @[Mux.scala 87:16]
  wire [31:0] op2_data; // @[Mux.scala 87:16]
  wire  _T_558; // @[Core.scala 163:52]
  wire  ecall_flg; // @[Core.scala 163:40]
  wire  _T_458; // @[Core.scala 132:18]
  wire [1:0] _T_189; // @[Lookup.scala 33:37]
  wire [1:0] _T_190; // @[Lookup.scala 33:37]
  wire [1:0] _T_191; // @[Lookup.scala 33:37]
  wire [1:0] _T_192; // @[Lookup.scala 33:37]
  wire [1:0] _T_193; // @[Lookup.scala 33:37]
  wire [1:0] _T_194; // @[Lookup.scala 33:37]
  wire [1:0] _T_195; // @[Lookup.scala 33:37]
  wire [1:0] _T_196; // @[Lookup.scala 33:37]
  wire [1:0] _T_197; // @[Lookup.scala 33:37]
  wire [1:0] _T_198; // @[Lookup.scala 33:37]
  wire [1:0] _T_199; // @[Lookup.scala 33:37]
  wire [1:0] _T_200; // @[Lookup.scala 33:37]
  wire [1:0] _T_201; // @[Lookup.scala 33:37]
  wire [1:0] _T_202; // @[Lookup.scala 33:37]
  wire [1:0] _T_203; // @[Lookup.scala 33:37]
  wire [1:0] _T_204; // @[Lookup.scala 33:37]
  wire [1:0] _T_205; // @[Lookup.scala 33:37]
  wire [1:0] _T_206; // @[Lookup.scala 33:37]
  wire [1:0] _T_207; // @[Lookup.scala 33:37]
  wire [1:0] _T_208; // @[Lookup.scala 33:37]
  wire [1:0] _T_209; // @[Lookup.scala 33:37]
  wire [1:0] _T_210; // @[Lookup.scala 33:37]
  wire [1:0] _T_211; // @[Lookup.scala 33:37]
  wire [1:0] _T_212; // @[Lookup.scala 33:37]
  wire [1:0] _T_213; // @[Lookup.scala 33:37]
  wire [1:0] _T_214; // @[Lookup.scala 33:37]
  wire [1:0] _T_215; // @[Lookup.scala 33:37]
  wire [1:0] _T_216; // @[Lookup.scala 33:37]
  wire [1:0] _T_217; // @[Lookup.scala 33:37]
  wire [1:0] _T_218; // @[Lookup.scala 33:37]
  wire [1:0] _T_219; // @[Lookup.scala 33:37]
  wire [1:0] _T_220; // @[Lookup.scala 33:37]
  wire [1:0] _T_221; // @[Lookup.scala 33:37]
  wire [1:0] _T_222; // @[Lookup.scala 33:37]
  wire [1:0] _T_223; // @[Lookup.scala 33:37]
  wire [1:0] _T_224; // @[Lookup.scala 33:37]
  wire [1:0] _T_225; // @[Lookup.scala 33:37]
  wire [1:0] _T_226; // @[Lookup.scala 33:37]
  wire [1:0] _T_227; // @[Lookup.scala 33:37]
  wire [1:0] _T_228; // @[Lookup.scala 33:37]
  wire [1:0] _T_229; // @[Lookup.scala 33:37]
  wire [1:0] _T_230; // @[Lookup.scala 33:37]
  wire [1:0] csignals_1; // @[Lookup.scala 33:37]
  wire  _T_446; // @[Core.scala 117:18]
  wire [4:0] rs1_addr; // @[Core.scala 40:24]
  wire  _T_15; // @[Core.scala 45:37]
  wire  _T_16; // @[Core.scala 45:25]
  wire [31:0] _T_17; // @[Mux.scala 87:16]
  wire [31:0] rs1_data; // @[Mux.scala 87:16]
  wire  _T_447; // @[Core.scala 118:18]
  wire [31:0] _T_448; // @[Mux.scala 87:16]
  wire [31:0] op1_data; // @[Mux.scala 87:16]
  wire [31:0] _T_460; // @[Core.scala 132:46]
  wire  _T_461; // @[Core.scala 133:18]
  wire [31:0] _T_463; // @[Core.scala 133:46]
  wire  _T_464; // @[Core.scala 134:18]
  wire [31:0] _T_465; // @[Core.scala 134:46]
  wire  _T_466; // @[Core.scala 135:18]
  wire [31:0] _T_467; // @[Core.scala 135:46]
  wire  _T_468; // @[Core.scala 136:18]
  wire [31:0] _T_469; // @[Core.scala 136:46]
  wire  _T_470; // @[Core.scala 137:18]
  wire [63:0] _T_471; // @[Core.scala 137:45]
  wire [31:0] _T_472; // @[Core.scala 137:56]
  wire  _T_473; // @[Core.scala 138:18]
  wire [31:0] _T_475; // @[Core.scala 138:55]
  wire  _T_476; // @[Core.scala 139:18]
  wire [31:0] _T_477; // @[Core.scala 139:50]
  wire [31:0] _T_478; // @[Core.scala 139:70]
  wire [32:0] _T_479; // @[Core.scala 139:53]
  wire [32:0] _T_480; // @[Core.scala 139:80]
  wire  _T_481; // @[Core.scala 140:18]
  wire [31:0] _T_482; // @[Core.scala 140:45]
  wire  _T_483; // @[Core.scala 141:18]
  wire [31:0] _GEN_0; // @[Core.scala 141:53]
  wire [31:0] _T_486; // @[Core.scala 141:53]
  wire [31:0] _T_487; // @[Core.scala 141:80]
  wire  _T_488; // @[Core.scala 142:18]
  wire [31:0] _GEN_1; // @[Core.scala 142:45]
  wire [31:0] _T_489; // @[Core.scala 142:45]
  wire  _T_490; // @[Core.scala 143:18]
  wire [4:0] _T_491; // @[Core.scala 143:57]
  wire [62:0] _GEN_5; // @[Core.scala 143:46]
  wire [62:0] _T_492; // @[Core.scala 143:46]
  wire [31:0] _T_493; // @[Core.scala 143:64]
  wire  _T_494; // @[Core.scala 144:18]
  wire [31:0] _T_496; // @[Core.scala 144:46]
  wire  _T_497; // @[Core.scala 145:18]
  wire [31:0] _T_500; // @[Core.scala 145:55]
  wire [31:0] _T_501; // @[Core.scala 145:80]
  wire  _T_502; // @[Core.scala 146:18]
  wire  _T_505; // @[Core.scala 146:55]
  wire  _T_506; // @[Core.scala 147:18]
  wire  _T_507; // @[Core.scala 147:46]
  wire  _T_508; // @[Core.scala 148:18]
  wire [31:0] _T_512; // @[Core.scala 148:59]
  wire [31:0] _T_513; // @[Mux.scala 87:16]
  wire [31:0] _T_514; // @[Mux.scala 87:16]
  wire [31:0] _T_515; // @[Mux.scala 87:16]
  wire [31:0] _T_516; // @[Mux.scala 87:16]
  wire [31:0] _T_517; // @[Mux.scala 87:16]
  wire [31:0] _T_518; // @[Mux.scala 87:16]
  wire [31:0] _T_519; // @[Mux.scala 87:16]
  wire [31:0] _T_520; // @[Mux.scala 87:16]
  wire [31:0] _T_521; // @[Mux.scala 87:16]
  wire [32:0] _T_522; // @[Mux.scala 87:16]
  wire [32:0] _T_523; // @[Mux.scala 87:16]
  wire [32:0] _T_524; // @[Mux.scala 87:16]
  wire [32:0] _T_525; // @[Mux.scala 87:16]
  wire [32:0] _T_526; // @[Mux.scala 87:16]
  wire [32:0] _T_527; // @[Mux.scala 87:16]
  wire [32:0] _T_528; // @[Mux.scala 87:16]
  wire [32:0] _T_529; // @[Mux.scala 87:16]
  wire [31:0] alu_out; // @[Core.scala 29:23 Core.scala 131:13]
  wire  _T_530; // @[Core.scala 153:18]
  wire  _T_531; // @[Core.scala 153:45]
  wire  _T_532; // @[Core.scala 154:18]
  wire  _T_534; // @[Core.scala 154:34]
  wire  _T_535; // @[Core.scala 155:18]
  wire  _T_539; // @[Core.scala 156:18]
  wire  _T_543; // @[Core.scala 156:34]
  wire  _T_544; // @[Core.scala 157:18]
  wire  _T_546; // @[Core.scala 158:18]
  wire  _T_548; // @[Core.scala 158:34]
  wire  _T_549; // @[Mux.scala 87:16]
  wire  _T_550; // @[Mux.scala 87:16]
  wire  _T_551; // @[Mux.scala 87:16]
  wire  _T_552; // @[Mux.scala 87:16]
  wire  _T_553; // @[Mux.scala 87:16]
  wire  br_flg; // @[Mux.scala 87:16]
  wire  _T_37; // @[Core.scala 57:35]
  wire [5:0] _T_38; // @[Core.scala 57:44]
  wire [3:0] _T_39; // @[Core.scala 57:58]
  wire [11:0] imm_b; // @[Cat.scala 29:58]
  wire  _T_42; // @[Core.scala 58:40]
  wire [18:0] _T_44; // @[Bitwise.scala 71:12]
  wire [31:0] imm_b_sext; // @[Cat.scala 29:58]
  wire [31:0] br_target; // @[Core.scala 160:25]
  wire [1:0] _T_310; // @[Lookup.scala 33:37]
  wire [1:0] _T_311; // @[Lookup.scala 33:37]
  wire [1:0] _T_312; // @[Lookup.scala 33:37]
  wire [1:0] _T_313; // @[Lookup.scala 33:37]
  wire [1:0] _T_314; // @[Lookup.scala 33:37]
  wire [1:0] _T_315; // @[Lookup.scala 33:37]
  wire [1:0] _T_316; // @[Lookup.scala 33:37]
  wire [1:0] csignals_3; // @[Lookup.scala 33:37]
  wire [1:0] _T_318; // @[Lookup.scala 33:37]
  wire [1:0] _T_319; // @[Lookup.scala 33:37]
  wire [1:0] _T_320; // @[Lookup.scala 33:37]
  wire [1:0] _T_321; // @[Lookup.scala 33:37]
  wire [1:0] _T_322; // @[Lookup.scala 33:37]
  wire [1:0] _T_323; // @[Lookup.scala 33:37]
  wire [1:0] _T_324; // @[Lookup.scala 33:37]
  wire [1:0] _T_325; // @[Lookup.scala 33:37]
  wire [1:0] _T_326; // @[Lookup.scala 33:37]
  wire [1:0] _T_327; // @[Lookup.scala 33:37]
  wire [1:0] _T_328; // @[Lookup.scala 33:37]
  wire [1:0] _T_329; // @[Lookup.scala 33:37]
  wire [1:0] _T_330; // @[Lookup.scala 33:37]
  wire [1:0] _T_331; // @[Lookup.scala 33:37]
  wire [1:0] _T_332; // @[Lookup.scala 33:37]
  wire [1:0] _T_333; // @[Lookup.scala 33:37]
  wire [1:0] _T_334; // @[Lookup.scala 33:37]
  wire [1:0] _T_335; // @[Lookup.scala 33:37]
  wire [1:0] _T_336; // @[Lookup.scala 33:37]
  wire [1:0] _T_337; // @[Lookup.scala 33:37]
  wire [1:0] _T_338; // @[Lookup.scala 33:37]
  wire [1:0] _T_339; // @[Lookup.scala 33:37]
  wire [1:0] _T_340; // @[Lookup.scala 33:37]
  wire [1:0] _T_341; // @[Lookup.scala 33:37]
  wire [1:0] _T_342; // @[Lookup.scala 33:37]
  wire [1:0] _T_343; // @[Lookup.scala 33:37]
  wire [1:0] _T_344; // @[Lookup.scala 33:37]
  wire [1:0] _T_345; // @[Lookup.scala 33:37]
  wire [1:0] _T_346; // @[Lookup.scala 33:37]
  wire [1:0] _T_347; // @[Lookup.scala 33:37]
  wire [1:0] _T_348; // @[Lookup.scala 33:37]
  wire [1:0] _T_349; // @[Lookup.scala 33:37]
  wire [1:0] _T_350; // @[Lookup.scala 33:37]
  wire [1:0] _T_351; // @[Lookup.scala 33:37]
  wire [1:0] _T_352; // @[Lookup.scala 33:37]
  wire [1:0] _T_353; // @[Lookup.scala 33:37]
  wire [1:0] _T_354; // @[Lookup.scala 33:37]
  wire [1:0] _T_355; // @[Lookup.scala 33:37]
  wire [1:0] _T_356; // @[Lookup.scala 33:37]
  wire [1:0] _T_357; // @[Lookup.scala 33:37]
  wire [1:0] _T_358; // @[Lookup.scala 33:37]
  wire [1:0] _T_359; // @[Lookup.scala 33:37]
  wire [1:0] csignals_4; // @[Lookup.scala 33:37]
  wire [2:0] _T_363; // @[Lookup.scala 33:37]
  wire [2:0] _T_364; // @[Lookup.scala 33:37]
  wire [2:0] _T_365; // @[Lookup.scala 33:37]
  wire [2:0] _T_366; // @[Lookup.scala 33:37]
  wire [2:0] _T_367; // @[Lookup.scala 33:37]
  wire [2:0] _T_368; // @[Lookup.scala 33:37]
  wire [2:0] _T_369; // @[Lookup.scala 33:37]
  wire [2:0] _T_370; // @[Lookup.scala 33:37]
  wire [2:0] _T_371; // @[Lookup.scala 33:37]
  wire [2:0] _T_372; // @[Lookup.scala 33:37]
  wire [2:0] _T_373; // @[Lookup.scala 33:37]
  wire [2:0] _T_374; // @[Lookup.scala 33:37]
  wire [2:0] _T_375; // @[Lookup.scala 33:37]
  wire [2:0] _T_376; // @[Lookup.scala 33:37]
  wire [2:0] _T_377; // @[Lookup.scala 33:37]
  wire [2:0] _T_378; // @[Lookup.scala 33:37]
  wire [2:0] _T_379; // @[Lookup.scala 33:37]
  wire [2:0] _T_380; // @[Lookup.scala 33:37]
  wire [2:0] _T_381; // @[Lookup.scala 33:37]
  wire [2:0] _T_382; // @[Lookup.scala 33:37]
  wire [2:0] _T_383; // @[Lookup.scala 33:37]
  wire [2:0] _T_384; // @[Lookup.scala 33:37]
  wire [2:0] _T_385; // @[Lookup.scala 33:37]
  wire [2:0] _T_386; // @[Lookup.scala 33:37]
  wire [2:0] _T_387; // @[Lookup.scala 33:37]
  wire [2:0] _T_388; // @[Lookup.scala 33:37]
  wire [2:0] _T_389; // @[Lookup.scala 33:37]
  wire [2:0] _T_390; // @[Lookup.scala 33:37]
  wire [2:0] _T_391; // @[Lookup.scala 33:37]
  wire [2:0] _T_392; // @[Lookup.scala 33:37]
  wire [2:0] _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_400; // @[Lookup.scala 33:37]
  wire [2:0] _T_401; // @[Lookup.scala 33:37]
  wire [2:0] _T_402; // @[Lookup.scala 33:37]
  wire [2:0] csignals_5; // @[Lookup.scala 33:37]
  wire [2:0] _T_439; // @[Lookup.scala 33:37]
  wire [2:0] _T_440; // @[Lookup.scala 33:37]
  wire [2:0] _T_441; // @[Lookup.scala 33:37]
  wire [2:0] _T_442; // @[Lookup.scala 33:37]
  wire [2:0] _T_443; // @[Lookup.scala 33:37]
  wire [2:0] _T_444; // @[Lookup.scala 33:37]
  wire [2:0] _T_445; // @[Lookup.scala 33:37]
  reg [31:0] seg_data; // @[Core.scala 164:27]
  reg [31:0] _RAND_2;
  wire  _T_561; // @[Core.scala 166:55]
  wire  _T_562; // @[Core.scala 166:43]
  wire  _T_564; // @[Core.scala 176:17]
  wire  _T_565; // @[Core.scala 177:17]
  wire [31:0] _T_566; // @[Mux.scala 87:16]
  assign regfile__T_8_addr = io_imem_inst[19:15];
  assign regfile__T_8_data = regfile[regfile__T_8_addr]; // @[Core.scala 17:22]
  assign regfile__T_11_addr = 5'ha;
  assign regfile__T_11_data = regfile[regfile__T_11_addr]; // @[Core.scala 17:22]
  assign regfile__T_18_addr = io_imem_inst[24:20];
  assign regfile__T_18_data = regfile[regfile__T_18_addr]; // @[Core.scala 17:22]
  assign regfile__T_21_addr = 5'h11;
  assign regfile__T_21_data = regfile[regfile__T_21_addr]; // @[Core.scala 17:22]
  assign regfile__T_568_data = _T_564 ? io_dmem_rdata : _T_566;
  assign regfile__T_568_addr = io_imem_inst[11:7];
  assign regfile__T_568_mask = 1'h1;
  assign regfile__T_568_en = csignals_4 == 2'h1;
  assign pc_plus4 = pc_reg + 32'h4; // @[Core.scala 25:27]
  assign _T_1 = io_imem_inst & 32'h7f; // @[Core.scala 33:15]
  assign _T_2 = 32'h6f == _T_1; // @[Core.scala 33:15]
  assign _T_3 = io_imem_inst & 32'h707f; // @[Core.scala 33:31]
  assign _T_4 = 32'h67 == _T_3; // @[Core.scala 33:31]
  assign _T_5 = _T_2 | _T_4; // @[Core.scala 33:23]
  assign _T_58 = 32'h3 == _T_3; // @[Lookup.scala 31:38]
  assign _T_60 = 32'h1003 == _T_3; // @[Lookup.scala 31:38]
  assign _T_62 = 32'h2003 == _T_3; // @[Lookup.scala 31:38]
  assign _T_64 = 32'h4003 == _T_3; // @[Lookup.scala 31:38]
  assign _T_66 = 32'h5003 == _T_3; // @[Lookup.scala 31:38]
  assign _T_68 = 32'h23 == _T_3; // @[Lookup.scala 31:38]
  assign _T_70 = 32'h1023 == _T_3; // @[Lookup.scala 31:38]
  assign _T_72 = 32'h2023 == _T_3; // @[Lookup.scala 31:38]
  assign _T_73 = io_imem_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  assign _T_74 = 32'h33 == _T_73; // @[Lookup.scala 31:38]
  assign _T_76 = 32'h13 == _T_3; // @[Lookup.scala 31:38]
  assign _T_78 = 32'h40000033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_80 = 32'h7033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_82 = 32'h6033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_84 = 32'h4033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_86 = 32'h7013 == _T_3; // @[Lookup.scala 31:38]
  assign _T_88 = 32'h6013 == _T_3; // @[Lookup.scala 31:38]
  assign _T_90 = 32'h4013 == _T_3; // @[Lookup.scala 31:38]
  assign _T_92 = 32'h2000033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_94 = 32'h2001033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_96 = 32'h2004033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_98 = 32'h2005033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_100 = 32'h2006033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_102 = 32'h2007033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_104 = 32'h1033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_106 = 32'h5033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_108 = 32'h40005033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_110 = 32'h1013 == _T_73; // @[Lookup.scala 31:38]
  assign _T_112 = 32'h5013 == _T_73; // @[Lookup.scala 31:38]
  assign _T_114 = 32'h40005013 == _T_73; // @[Lookup.scala 31:38]
  assign _T_116 = 32'h2033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_118 = 32'h3033 == _T_73; // @[Lookup.scala 31:38]
  assign _T_120 = 32'h2013 == _T_3; // @[Lookup.scala 31:38]
  assign _T_122 = 32'h3013 == _T_3; // @[Lookup.scala 31:38]
  assign _T_124 = 32'h63 == _T_3; // @[Lookup.scala 31:38]
  assign _T_126 = 32'h1063 == _T_3; // @[Lookup.scala 31:38]
  assign _T_128 = 32'h5063 == _T_3; // @[Lookup.scala 31:38]
  assign _T_130 = 32'h7063 == _T_3; // @[Lookup.scala 31:38]
  assign _T_132 = 32'h4063 == _T_3; // @[Lookup.scala 31:38]
  assign _T_134 = 32'h6063 == _T_3; // @[Lookup.scala 31:38]
  assign _T_140 = 32'h37 == _T_1; // @[Lookup.scala 31:38]
  assign _T_142 = 32'h17 == _T_1; // @[Lookup.scala 31:38]
  assign _T_144 = 32'h73 == io_imem_inst; // @[Lookup.scala 31:38]
  assign _T_145 = _T_144 ? 5'h18 : 5'h0; // @[Lookup.scala 33:37]
  assign _T_146 = _T_142 ? 5'h1 : _T_145; // @[Lookup.scala 33:37]
  assign _T_147 = _T_140 ? 5'h1 : _T_146; // @[Lookup.scala 33:37]
  assign _T_148 = _T_4 ? 5'h11 : _T_147; // @[Lookup.scala 33:37]
  assign _T_149 = _T_2 ? 5'h1 : _T_148; // @[Lookup.scala 33:37]
  assign _T_150 = _T_134 ? 5'hf : _T_149; // @[Lookup.scala 33:37]
  assign _T_151 = _T_132 ? 5'hd : _T_150; // @[Lookup.scala 33:37]
  assign _T_152 = _T_130 ? 5'h10 : _T_151; // @[Lookup.scala 33:37]
  assign _T_153 = _T_128 ? 5'he : _T_152; // @[Lookup.scala 33:37]
  assign _T_154 = _T_126 ? 5'hc : _T_153; // @[Lookup.scala 33:37]
  assign _T_155 = _T_124 ? 5'hb : _T_154; // @[Lookup.scala 33:37]
  assign _T_156 = _T_122 ? 5'ha : _T_155; // @[Lookup.scala 33:37]
  assign _T_157 = _T_120 ? 5'h9 : _T_156; // @[Lookup.scala 33:37]
  assign _T_158 = _T_118 ? 5'ha : _T_157; // @[Lookup.scala 33:37]
  assign _T_159 = _T_116 ? 5'h9 : _T_158; // @[Lookup.scala 33:37]
  assign _T_160 = _T_114 ? 5'h8 : _T_159; // @[Lookup.scala 33:37]
  assign _T_161 = _T_112 ? 5'h7 : _T_160; // @[Lookup.scala 33:37]
  assign _T_162 = _T_110 ? 5'h6 : _T_161; // @[Lookup.scala 33:37]
  assign _T_163 = _T_108 ? 5'h8 : _T_162; // @[Lookup.scala 33:37]
  assign _T_164 = _T_106 ? 5'h7 : _T_163; // @[Lookup.scala 33:37]
  assign _T_165 = _T_104 ? 5'h6 : _T_164; // @[Lookup.scala 33:37]
  assign _T_166 = _T_102 ? 5'h17 : _T_165; // @[Lookup.scala 33:37]
  assign _T_167 = _T_100 ? 5'h16 : _T_166; // @[Lookup.scala 33:37]
  assign _T_168 = _T_98 ? 5'h15 : _T_167; // @[Lookup.scala 33:37]
  assign _T_169 = _T_96 ? 5'h14 : _T_168; // @[Lookup.scala 33:37]
  assign _T_170 = _T_94 ? 5'h13 : _T_169; // @[Lookup.scala 33:37]
  assign _T_171 = _T_92 ? 5'h12 : _T_170; // @[Lookup.scala 33:37]
  assign _T_172 = _T_90 ? 5'h5 : _T_171; // @[Lookup.scala 33:37]
  assign _T_173 = _T_88 ? 5'h4 : _T_172; // @[Lookup.scala 33:37]
  assign _T_174 = _T_86 ? 5'h3 : _T_173; // @[Lookup.scala 33:37]
  assign _T_175 = _T_84 ? 5'h5 : _T_174; // @[Lookup.scala 33:37]
  assign _T_176 = _T_82 ? 5'h4 : _T_175; // @[Lookup.scala 33:37]
  assign _T_177 = _T_80 ? 5'h3 : _T_176; // @[Lookup.scala 33:37]
  assign _T_178 = _T_78 ? 5'h2 : _T_177; // @[Lookup.scala 33:37]
  assign _T_179 = _T_76 ? 5'h1 : _T_178; // @[Lookup.scala 33:37]
  assign _T_180 = _T_74 ? 5'h1 : _T_179; // @[Lookup.scala 33:37]
  assign _T_181 = _T_72 ? 5'h1 : _T_180; // @[Lookup.scala 33:37]
  assign _T_182 = _T_70 ? 5'h1 : _T_181; // @[Lookup.scala 33:37]
  assign _T_183 = _T_68 ? 5'h1 : _T_182; // @[Lookup.scala 33:37]
  assign _T_184 = _T_66 ? 5'h1 : _T_183; // @[Lookup.scala 33:37]
  assign _T_185 = _T_64 ? 5'h1 : _T_184; // @[Lookup.scala 33:37]
  assign _T_186 = _T_62 ? 5'h1 : _T_185; // @[Lookup.scala 33:37]
  assign _T_187 = _T_60 ? 5'h1 : _T_186; // @[Lookup.scala 33:37]
  assign csignals_0 = _T_58 ? 5'h1 : _T_187; // @[Lookup.scala 33:37]
  assign _T_557 = csignals_0 == 5'h18; // @[Core.scala 163:27]
  assign _T_232 = _T_142 ? 3'h5 : 3'h1; // @[Lookup.scala 33:37]
  assign _T_233 = _T_140 ? 3'h5 : _T_232; // @[Lookup.scala 33:37]
  assign _T_234 = _T_4 ? 3'h2 : _T_233; // @[Lookup.scala 33:37]
  assign _T_235 = _T_2 ? 3'h4 : _T_234; // @[Lookup.scala 33:37]
  assign _T_236 = _T_134 ? 3'h1 : _T_235; // @[Lookup.scala 33:37]
  assign _T_237 = _T_132 ? 3'h1 : _T_236; // @[Lookup.scala 33:37]
  assign _T_238 = _T_130 ? 3'h1 : _T_237; // @[Lookup.scala 33:37]
  assign _T_239 = _T_128 ? 3'h1 : _T_238; // @[Lookup.scala 33:37]
  assign _T_240 = _T_126 ? 3'h1 : _T_239; // @[Lookup.scala 33:37]
  assign _T_241 = _T_124 ? 3'h1 : _T_240; // @[Lookup.scala 33:37]
  assign _T_242 = _T_122 ? 3'h2 : _T_241; // @[Lookup.scala 33:37]
  assign _T_243 = _T_120 ? 3'h2 : _T_242; // @[Lookup.scala 33:37]
  assign _T_244 = _T_118 ? 3'h1 : _T_243; // @[Lookup.scala 33:37]
  assign _T_245 = _T_116 ? 3'h1 : _T_244; // @[Lookup.scala 33:37]
  assign _T_246 = _T_114 ? 3'h2 : _T_245; // @[Lookup.scala 33:37]
  assign _T_247 = _T_112 ? 3'h2 : _T_246; // @[Lookup.scala 33:37]
  assign _T_248 = _T_110 ? 3'h2 : _T_247; // @[Lookup.scala 33:37]
  assign _T_249 = _T_108 ? 3'h1 : _T_248; // @[Lookup.scala 33:37]
  assign _T_250 = _T_106 ? 3'h1 : _T_249; // @[Lookup.scala 33:37]
  assign _T_251 = _T_104 ? 3'h1 : _T_250; // @[Lookup.scala 33:37]
  assign _T_252 = _T_102 ? 3'h1 : _T_251; // @[Lookup.scala 33:37]
  assign _T_253 = _T_100 ? 3'h1 : _T_252; // @[Lookup.scala 33:37]
  assign _T_254 = _T_98 ? 3'h1 : _T_253; // @[Lookup.scala 33:37]
  assign _T_255 = _T_96 ? 3'h1 : _T_254; // @[Lookup.scala 33:37]
  assign _T_256 = _T_94 ? 3'h1 : _T_255; // @[Lookup.scala 33:37]
  assign _T_257 = _T_92 ? 3'h1 : _T_256; // @[Lookup.scala 33:37]
  assign _T_258 = _T_90 ? 3'h2 : _T_257; // @[Lookup.scala 33:37]
  assign _T_259 = _T_88 ? 3'h2 : _T_258; // @[Lookup.scala 33:37]
  assign _T_260 = _T_86 ? 3'h2 : _T_259; // @[Lookup.scala 33:37]
  assign _T_261 = _T_84 ? 3'h1 : _T_260; // @[Lookup.scala 33:37]
  assign _T_262 = _T_82 ? 3'h1 : _T_261; // @[Lookup.scala 33:37]
  assign _T_263 = _T_80 ? 3'h1 : _T_262; // @[Lookup.scala 33:37]
  assign _T_264 = _T_78 ? 3'h1 : _T_263; // @[Lookup.scala 33:37]
  assign _T_265 = _T_76 ? 3'h2 : _T_264; // @[Lookup.scala 33:37]
  assign _T_266 = _T_74 ? 3'h1 : _T_265; // @[Lookup.scala 33:37]
  assign _T_267 = _T_72 ? 3'h3 : _T_266; // @[Lookup.scala 33:37]
  assign _T_268 = _T_70 ? 3'h3 : _T_267; // @[Lookup.scala 33:37]
  assign _T_269 = _T_68 ? 3'h3 : _T_268; // @[Lookup.scala 33:37]
  assign _T_270 = _T_66 ? 3'h2 : _T_269; // @[Lookup.scala 33:37]
  assign _T_271 = _T_64 ? 3'h2 : _T_270; // @[Lookup.scala 33:37]
  assign _T_272 = _T_62 ? 3'h2 : _T_271; // @[Lookup.scala 33:37]
  assign _T_273 = _T_60 ? 3'h2 : _T_272; // @[Lookup.scala 33:37]
  assign csignals_2 = _T_58 ? 3'h2 : _T_273; // @[Lookup.scala 33:37]
  assign _T_449 = csignals_2 == 3'h1; // @[Core.scala 122:18]
  assign _T_24 = _T_144 == 1'h0; // @[Core.scala 50:15]
  assign rs2_addr = io_imem_inst[24:20]; // @[Core.scala 41:24]
  assign _T_25 = rs2_addr == 5'h0; // @[Core.scala 50:37]
  assign _T_26 = _T_24 & _T_25; // @[Core.scala 50:25]
  assign _T_27 = _T_26 ? 32'h0 : regfile__T_18_data; // @[Mux.scala 87:16]
  assign rs2_data = _T_144 ? regfile__T_21_data : _T_27; // @[Mux.scala 87:16]
  assign _T_450 = csignals_2 == 3'h2; // @[Core.scala 123:18]
  assign imm_i = io_imem_inst[31:20]; // @[Core.scala 53:21]
  assign _T_28 = imm_i[11]; // @[Core.scala 54:40]
  assign _T_30 = _T_28 ? 20'hfffff : 20'h0; // @[Bitwise.scala 71:12]
  assign imm_i_sext = {_T_30,imm_i}; // @[Cat.scala 29:58]
  assign _T_451 = csignals_2 == 3'h3; // @[Core.scala 124:18]
  assign _T_31 = io_imem_inst[31:25]; // @[Core.scala 55:25]
  assign _T_32 = io_imem_inst[11:7]; // @[Core.scala 55:39]
  assign imm_s = {_T_31,_T_32}; // @[Cat.scala 29:58]
  assign _T_33 = imm_s[11]; // @[Core.scala 56:40]
  assign _T_35 = _T_33 ? 20'hfffff : 20'h0; // @[Bitwise.scala 71:12]
  assign imm_s_sext = {_T_35,_T_31,_T_32}; // @[Cat.scala 29:58]
  assign _T_452 = csignals_2 == 3'h4; // @[Core.scala 125:18]
  assign _T_46 = io_imem_inst[31]; // @[Core.scala 59:25]
  assign _T_47 = io_imem_inst[19:12]; // @[Core.scala 59:35]
  assign _T_48 = io_imem_inst[20]; // @[Core.scala 59:49]
  assign _T_49 = io_imem_inst[30:21]; // @[Core.scala 59:59]
  assign imm_j = {_T_46,_T_47,_T_48,_T_49}; // @[Cat.scala 29:58]
  assign _T_52 = imm_j[19]; // @[Core.scala 60:40]
  assign _T_54 = _T_52 ? 11'h7ff : 11'h0; // @[Bitwise.scala 71:12]
  assign imm_j_sext = {_T_54,_T_46,_T_47,_T_48,_T_49,1'h0}; // @[Cat.scala 29:58]
  assign _T_453 = csignals_2 == 3'h5; // @[Core.scala 126:18]
  assign imm_u = io_imem_inst[31:12]; // @[Core.scala 61:21]
  assign imm_u_shifted = {imm_u,12'h0}; // @[Cat.scala 29:58]
  assign _T_454 = _T_453 ? imm_u_shifted : 32'h0; // @[Mux.scala 87:16]
  assign _T_455 = _T_452 ? imm_j_sext : _T_454; // @[Mux.scala 87:16]
  assign _T_456 = _T_451 ? imm_s_sext : _T_455; // @[Mux.scala 87:16]
  assign _T_457 = _T_450 ? imm_i_sext : _T_456; // @[Mux.scala 87:16]
  assign op2_data = _T_449 ? rs2_data : _T_457; // @[Mux.scala 87:16]
  assign _T_558 = op2_data != 32'h22; // @[Core.scala 163:52]
  assign ecall_flg = _T_557 & _T_558; // @[Core.scala 163:40]
  assign _T_458 = csignals_0 == 5'h1; // @[Core.scala 132:18]
  assign _T_189 = _T_142 ? 2'h2 : 2'h1; // @[Lookup.scala 33:37]
  assign _T_190 = _T_140 ? 2'h0 : _T_189; // @[Lookup.scala 33:37]
  assign _T_191 = _T_4 ? 2'h1 : _T_190; // @[Lookup.scala 33:37]
  assign _T_192 = _T_2 ? 2'h2 : _T_191; // @[Lookup.scala 33:37]
  assign _T_193 = _T_134 ? 2'h1 : _T_192; // @[Lookup.scala 33:37]
  assign _T_194 = _T_132 ? 2'h1 : _T_193; // @[Lookup.scala 33:37]
  assign _T_195 = _T_130 ? 2'h1 : _T_194; // @[Lookup.scala 33:37]
  assign _T_196 = _T_128 ? 2'h1 : _T_195; // @[Lookup.scala 33:37]
  assign _T_197 = _T_126 ? 2'h1 : _T_196; // @[Lookup.scala 33:37]
  assign _T_198 = _T_124 ? 2'h1 : _T_197; // @[Lookup.scala 33:37]
  assign _T_199 = _T_122 ? 2'h1 : _T_198; // @[Lookup.scala 33:37]
  assign _T_200 = _T_120 ? 2'h1 : _T_199; // @[Lookup.scala 33:37]
  assign _T_201 = _T_118 ? 2'h1 : _T_200; // @[Lookup.scala 33:37]
  assign _T_202 = _T_116 ? 2'h1 : _T_201; // @[Lookup.scala 33:37]
  assign _T_203 = _T_114 ? 2'h1 : _T_202; // @[Lookup.scala 33:37]
  assign _T_204 = _T_112 ? 2'h1 : _T_203; // @[Lookup.scala 33:37]
  assign _T_205 = _T_110 ? 2'h1 : _T_204; // @[Lookup.scala 33:37]
  assign _T_206 = _T_108 ? 2'h1 : _T_205; // @[Lookup.scala 33:37]
  assign _T_207 = _T_106 ? 2'h1 : _T_206; // @[Lookup.scala 33:37]
  assign _T_208 = _T_104 ? 2'h1 : _T_207; // @[Lookup.scala 33:37]
  assign _T_209 = _T_102 ? 2'h1 : _T_208; // @[Lookup.scala 33:37]
  assign _T_210 = _T_100 ? 2'h1 : _T_209; // @[Lookup.scala 33:37]
  assign _T_211 = _T_98 ? 2'h1 : _T_210; // @[Lookup.scala 33:37]
  assign _T_212 = _T_96 ? 2'h1 : _T_211; // @[Lookup.scala 33:37]
  assign _T_213 = _T_94 ? 2'h1 : _T_212; // @[Lookup.scala 33:37]
  assign _T_214 = _T_92 ? 2'h1 : _T_213; // @[Lookup.scala 33:37]
  assign _T_215 = _T_90 ? 2'h1 : _T_214; // @[Lookup.scala 33:37]
  assign _T_216 = _T_88 ? 2'h1 : _T_215; // @[Lookup.scala 33:37]
  assign _T_217 = _T_86 ? 2'h1 : _T_216; // @[Lookup.scala 33:37]
  assign _T_218 = _T_84 ? 2'h1 : _T_217; // @[Lookup.scala 33:37]
  assign _T_219 = _T_82 ? 2'h1 : _T_218; // @[Lookup.scala 33:37]
  assign _T_220 = _T_80 ? 2'h1 : _T_219; // @[Lookup.scala 33:37]
  assign _T_221 = _T_78 ? 2'h1 : _T_220; // @[Lookup.scala 33:37]
  assign _T_222 = _T_76 ? 2'h1 : _T_221; // @[Lookup.scala 33:37]
  assign _T_223 = _T_74 ? 2'h1 : _T_222; // @[Lookup.scala 33:37]
  assign _T_224 = _T_72 ? 2'h1 : _T_223; // @[Lookup.scala 33:37]
  assign _T_225 = _T_70 ? 2'h1 : _T_224; // @[Lookup.scala 33:37]
  assign _T_226 = _T_68 ? 2'h1 : _T_225; // @[Lookup.scala 33:37]
  assign _T_227 = _T_66 ? 2'h1 : _T_226; // @[Lookup.scala 33:37]
  assign _T_228 = _T_64 ? 2'h1 : _T_227; // @[Lookup.scala 33:37]
  assign _T_229 = _T_62 ? 2'h1 : _T_228; // @[Lookup.scala 33:37]
  assign _T_230 = _T_60 ? 2'h1 : _T_229; // @[Lookup.scala 33:37]
  assign csignals_1 = _T_58 ? 2'h1 : _T_230; // @[Lookup.scala 33:37]
  assign _T_446 = csignals_1 == 2'h1; // @[Core.scala 117:18]
  assign rs1_addr = io_imem_inst[19:15]; // @[Core.scala 40:24]
  assign _T_15 = rs1_addr == 5'h0; // @[Core.scala 45:37]
  assign _T_16 = _T_24 & _T_15; // @[Core.scala 45:25]
  assign _T_17 = _T_16 ? 32'h0 : regfile__T_8_data; // @[Mux.scala 87:16]
  assign rs1_data = _T_144 ? regfile__T_11_data : _T_17; // @[Mux.scala 87:16]
  assign _T_447 = csignals_1 == 2'h2; // @[Core.scala 118:18]
  assign _T_448 = _T_447 ? pc_reg : 32'h0; // @[Mux.scala 87:16]
  assign op1_data = _T_446 ? rs1_data : _T_448; // @[Mux.scala 87:16]
  assign _T_460 = op1_data + op2_data; // @[Core.scala 132:46]
  assign _T_461 = csignals_0 == 5'h2; // @[Core.scala 133:18]
  assign _T_463 = op1_data - op2_data; // @[Core.scala 133:46]
  assign _T_464 = csignals_0 == 5'h3; // @[Core.scala 134:18]
  assign _T_465 = op1_data & op2_data; // @[Core.scala 134:46]
  assign _T_466 = csignals_0 == 5'h4; // @[Core.scala 135:18]
  assign _T_467 = op1_data | op2_data; // @[Core.scala 135:46]
  assign _T_468 = csignals_0 == 5'h5; // @[Core.scala 136:18]
  assign _T_469 = op1_data ^ op2_data; // @[Core.scala 136:46]
  assign _T_470 = csignals_0 == 5'h12; // @[Core.scala 137:18]
  assign _T_471 = op1_data * op2_data; // @[Core.scala 137:45]
  assign _T_472 = _T_471[31:0]; // @[Core.scala 137:56]
  assign _T_473 = csignals_0 == 5'h13; // @[Core.scala 138:18]
  assign _T_475 = _T_471[63:32]; // @[Core.scala 138:55]
  assign _T_476 = csignals_0 == 5'h14; // @[Core.scala 139:18]
  assign _T_477 = $signed(op1_data); // @[Core.scala 139:50]
  assign _T_478 = $signed(op2_data); // @[Core.scala 139:70]
  assign _T_479 = $signed(_T_477) / $signed(_T_478); // @[Core.scala 139:53]
  assign _T_480 = $unsigned(_T_479); // @[Core.scala 139:80]
  assign _T_481 = csignals_0 == 5'h15; // @[Core.scala 140:18]
  assign _T_482 = op1_data / op2_data; // @[Core.scala 140:45]
  assign _T_483 = csignals_0 == 5'h16; // @[Core.scala 141:18]
  assign _GEN_0 = $signed(_T_477) % $signed(_T_478); // @[Core.scala 141:53]
  assign _T_486 = _GEN_0[31:0]; // @[Core.scala 141:53]
  assign _T_487 = $unsigned(_T_486); // @[Core.scala 141:80]
  assign _T_488 = csignals_0 == 5'h17; // @[Core.scala 142:18]
  assign _GEN_1 = op1_data % op2_data; // @[Core.scala 142:45]
  assign _T_489 = _GEN_1[31:0]; // @[Core.scala 142:45]
  assign _T_490 = csignals_0 == 5'h6; // @[Core.scala 143:18]
  assign _T_491 = op2_data[4:0]; // @[Core.scala 143:57]
  assign _GEN_5 = {{31'd0}, op1_data}; // @[Core.scala 143:46]
  assign _T_492 = _GEN_5 << _T_491; // @[Core.scala 143:46]
  assign _T_493 = _T_492[31:0]; // @[Core.scala 143:64]
  assign _T_494 = csignals_0 == 5'h7; // @[Core.scala 144:18]
  assign _T_496 = op1_data >> _T_491; // @[Core.scala 144:46]
  assign _T_497 = csignals_0 == 5'h8; // @[Core.scala 145:18]
  assign _T_500 = $signed(_T_477) >>> _T_491; // @[Core.scala 145:55]
  assign _T_501 = $unsigned(_T_500); // @[Core.scala 145:80]
  assign _T_502 = csignals_0 == 5'h9; // @[Core.scala 146:18]
  assign _T_505 = $signed(_T_477) < $signed(_T_478); // @[Core.scala 146:55]
  assign _T_506 = csignals_0 == 5'ha; // @[Core.scala 147:18]
  assign _T_507 = op1_data < op2_data; // @[Core.scala 147:46]
  assign _T_508 = csignals_0 == 5'h11; // @[Core.scala 148:18]
  assign _T_512 = _T_460 & 32'hfffffffe; // @[Core.scala 148:59]
  assign _T_513 = _T_508 ? _T_512 : 32'h0; // @[Mux.scala 87:16]
  assign _T_514 = _T_506 ? {{31'd0}, _T_507} : _T_513; // @[Mux.scala 87:16]
  assign _T_515 = _T_502 ? {{31'd0}, _T_505} : _T_514; // @[Mux.scala 87:16]
  assign _T_516 = _T_497 ? _T_501 : _T_515; // @[Mux.scala 87:16]
  assign _T_517 = _T_494 ? _T_496 : _T_516; // @[Mux.scala 87:16]
  assign _T_518 = _T_490 ? _T_493 : _T_517; // @[Mux.scala 87:16]
  assign _T_519 = _T_488 ? _T_489 : _T_518; // @[Mux.scala 87:16]
  assign _T_520 = _T_483 ? _T_487 : _T_519; // @[Mux.scala 87:16]
  assign _T_521 = _T_481 ? _T_482 : _T_520; // @[Mux.scala 87:16]
  assign _T_522 = _T_476 ? _T_480 : {{1'd0}, _T_521}; // @[Mux.scala 87:16]
  assign _T_523 = _T_473 ? {{1'd0}, _T_475} : _T_522; // @[Mux.scala 87:16]
  assign _T_524 = _T_470 ? {{1'd0}, _T_472} : _T_523; // @[Mux.scala 87:16]
  assign _T_525 = _T_468 ? {{1'd0}, _T_469} : _T_524; // @[Mux.scala 87:16]
  assign _T_526 = _T_466 ? {{1'd0}, _T_467} : _T_525; // @[Mux.scala 87:16]
  assign _T_527 = _T_464 ? {{1'd0}, _T_465} : _T_526; // @[Mux.scala 87:16]
  assign _T_528 = _T_461 ? {{1'd0}, _T_463} : _T_527; // @[Mux.scala 87:16]
  assign _T_529 = _T_458 ? {{1'd0}, _T_460} : _T_528; // @[Mux.scala 87:16]
  assign alu_out = _T_529[31:0]; // @[Core.scala 29:23 Core.scala 131:13]
  assign _T_530 = csignals_0 == 5'hb; // @[Core.scala 153:18]
  assign _T_531 = op1_data == op2_data; // @[Core.scala 153:45]
  assign _T_532 = csignals_0 == 5'hc; // @[Core.scala 154:18]
  assign _T_534 = _T_531 == 1'h0; // @[Core.scala 154:34]
  assign _T_535 = csignals_0 == 5'hd; // @[Core.scala 155:18]
  assign _T_539 = csignals_0 == 5'he; // @[Core.scala 156:18]
  assign _T_543 = _T_505 == 1'h0; // @[Core.scala 156:34]
  assign _T_544 = csignals_0 == 5'hf; // @[Core.scala 157:18]
  assign _T_546 = csignals_0 == 5'h10; // @[Core.scala 158:18]
  assign _T_548 = _T_507 == 1'h0; // @[Core.scala 158:34]
  assign _T_549 = _T_546 & _T_548; // @[Mux.scala 87:16]
  assign _T_550 = _T_544 ? _T_507 : _T_549; // @[Mux.scala 87:16]
  assign _T_551 = _T_539 ? _T_543 : _T_550; // @[Mux.scala 87:16]
  assign _T_552 = _T_535 ? _T_505 : _T_551; // @[Mux.scala 87:16]
  assign _T_553 = _T_532 ? _T_534 : _T_552; // @[Mux.scala 87:16]
  assign br_flg = _T_530 ? _T_531 : _T_553; // @[Mux.scala 87:16]
  assign _T_37 = io_imem_inst[7]; // @[Core.scala 57:35]
  assign _T_38 = io_imem_inst[30:25]; // @[Core.scala 57:44]
  assign _T_39 = io_imem_inst[11:8]; // @[Core.scala 57:58]
  assign imm_b = {_T_46,_T_37,_T_38,_T_39}; // @[Cat.scala 29:58]
  assign _T_42 = imm_b[11]; // @[Core.scala 58:40]
  assign _T_44 = _T_42 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 71:12]
  assign imm_b_sext = {_T_44,_T_46,_T_37,_T_38,_T_39,1'h0}; // @[Cat.scala 29:58]
  assign br_target = pc_reg + imm_b_sext; // @[Core.scala 160:25]
  assign _T_310 = _T_72 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  assign _T_311 = _T_70 ? 2'h1 : _T_310; // @[Lookup.scala 33:37]
  assign _T_312 = _T_68 ? 2'h1 : _T_311; // @[Lookup.scala 33:37]
  assign _T_313 = _T_66 ? 2'h0 : _T_312; // @[Lookup.scala 33:37]
  assign _T_314 = _T_64 ? 2'h0 : _T_313; // @[Lookup.scala 33:37]
  assign _T_315 = _T_62 ? 2'h0 : _T_314; // @[Lookup.scala 33:37]
  assign _T_316 = _T_60 ? 2'h0 : _T_315; // @[Lookup.scala 33:37]
  assign csignals_3 = _T_58 ? 2'h0 : _T_316; // @[Lookup.scala 33:37]
  assign _T_318 = _T_142 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  assign _T_319 = _T_140 ? 2'h1 : _T_318; // @[Lookup.scala 33:37]
  assign _T_320 = _T_4 ? 2'h1 : _T_319; // @[Lookup.scala 33:37]
  assign _T_321 = _T_2 ? 2'h1 : _T_320; // @[Lookup.scala 33:37]
  assign _T_322 = _T_134 ? 2'h0 : _T_321; // @[Lookup.scala 33:37]
  assign _T_323 = _T_132 ? 2'h0 : _T_322; // @[Lookup.scala 33:37]
  assign _T_324 = _T_130 ? 2'h0 : _T_323; // @[Lookup.scala 33:37]
  assign _T_325 = _T_128 ? 2'h0 : _T_324; // @[Lookup.scala 33:37]
  assign _T_326 = _T_126 ? 2'h0 : _T_325; // @[Lookup.scala 33:37]
  assign _T_327 = _T_124 ? 2'h0 : _T_326; // @[Lookup.scala 33:37]
  assign _T_328 = _T_122 ? 2'h1 : _T_327; // @[Lookup.scala 33:37]
  assign _T_329 = _T_120 ? 2'h1 : _T_328; // @[Lookup.scala 33:37]
  assign _T_330 = _T_118 ? 2'h1 : _T_329; // @[Lookup.scala 33:37]
  assign _T_331 = _T_116 ? 2'h1 : _T_330; // @[Lookup.scala 33:37]
  assign _T_332 = _T_114 ? 2'h1 : _T_331; // @[Lookup.scala 33:37]
  assign _T_333 = _T_112 ? 2'h1 : _T_332; // @[Lookup.scala 33:37]
  assign _T_334 = _T_110 ? 2'h1 : _T_333; // @[Lookup.scala 33:37]
  assign _T_335 = _T_108 ? 2'h1 : _T_334; // @[Lookup.scala 33:37]
  assign _T_336 = _T_106 ? 2'h1 : _T_335; // @[Lookup.scala 33:37]
  assign _T_337 = _T_104 ? 2'h1 : _T_336; // @[Lookup.scala 33:37]
  assign _T_338 = _T_102 ? 2'h1 : _T_337; // @[Lookup.scala 33:37]
  assign _T_339 = _T_100 ? 2'h1 : _T_338; // @[Lookup.scala 33:37]
  assign _T_340 = _T_98 ? 2'h1 : _T_339; // @[Lookup.scala 33:37]
  assign _T_341 = _T_96 ? 2'h1 : _T_340; // @[Lookup.scala 33:37]
  assign _T_342 = _T_94 ? 2'h1 : _T_341; // @[Lookup.scala 33:37]
  assign _T_343 = _T_92 ? 2'h1 : _T_342; // @[Lookup.scala 33:37]
  assign _T_344 = _T_90 ? 2'h1 : _T_343; // @[Lookup.scala 33:37]
  assign _T_345 = _T_88 ? 2'h1 : _T_344; // @[Lookup.scala 33:37]
  assign _T_346 = _T_86 ? 2'h1 : _T_345; // @[Lookup.scala 33:37]
  assign _T_347 = _T_84 ? 2'h1 : _T_346; // @[Lookup.scala 33:37]
  assign _T_348 = _T_82 ? 2'h1 : _T_347; // @[Lookup.scala 33:37]
  assign _T_349 = _T_80 ? 2'h1 : _T_348; // @[Lookup.scala 33:37]
  assign _T_350 = _T_78 ? 2'h1 : _T_349; // @[Lookup.scala 33:37]
  assign _T_351 = _T_76 ? 2'h1 : _T_350; // @[Lookup.scala 33:37]
  assign _T_352 = _T_74 ? 2'h1 : _T_351; // @[Lookup.scala 33:37]
  assign _T_353 = _T_72 ? 2'h0 : _T_352; // @[Lookup.scala 33:37]
  assign _T_354 = _T_70 ? 2'h0 : _T_353; // @[Lookup.scala 33:37]
  assign _T_355 = _T_68 ? 2'h0 : _T_354; // @[Lookup.scala 33:37]
  assign _T_356 = _T_66 ? 2'h1 : _T_355; // @[Lookup.scala 33:37]
  assign _T_357 = _T_64 ? 2'h1 : _T_356; // @[Lookup.scala 33:37]
  assign _T_358 = _T_62 ? 2'h1 : _T_357; // @[Lookup.scala 33:37]
  assign _T_359 = _T_60 ? 2'h1 : _T_358; // @[Lookup.scala 33:37]
  assign csignals_4 = _T_58 ? 2'h1 : _T_359; // @[Lookup.scala 33:37]
  assign _T_363 = _T_4 ? 3'h2 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_364 = _T_2 ? 3'h2 : _T_363; // @[Lookup.scala 33:37]
  assign _T_365 = _T_134 ? 3'h0 : _T_364; // @[Lookup.scala 33:37]
  assign _T_366 = _T_132 ? 3'h0 : _T_365; // @[Lookup.scala 33:37]
  assign _T_367 = _T_130 ? 3'h0 : _T_366; // @[Lookup.scala 33:37]
  assign _T_368 = _T_128 ? 3'h0 : _T_367; // @[Lookup.scala 33:37]
  assign _T_369 = _T_126 ? 3'h0 : _T_368; // @[Lookup.scala 33:37]
  assign _T_370 = _T_124 ? 3'h0 : _T_369; // @[Lookup.scala 33:37]
  assign _T_371 = _T_122 ? 3'h0 : _T_370; // @[Lookup.scala 33:37]
  assign _T_372 = _T_120 ? 3'h0 : _T_371; // @[Lookup.scala 33:37]
  assign _T_373 = _T_118 ? 3'h0 : _T_372; // @[Lookup.scala 33:37]
  assign _T_374 = _T_116 ? 3'h0 : _T_373; // @[Lookup.scala 33:37]
  assign _T_375 = _T_114 ? 3'h0 : _T_374; // @[Lookup.scala 33:37]
  assign _T_376 = _T_112 ? 3'h0 : _T_375; // @[Lookup.scala 33:37]
  assign _T_377 = _T_110 ? 3'h0 : _T_376; // @[Lookup.scala 33:37]
  assign _T_378 = _T_108 ? 3'h0 : _T_377; // @[Lookup.scala 33:37]
  assign _T_379 = _T_106 ? 3'h0 : _T_378; // @[Lookup.scala 33:37]
  assign _T_380 = _T_104 ? 3'h0 : _T_379; // @[Lookup.scala 33:37]
  assign _T_381 = _T_102 ? 3'h0 : _T_380; // @[Lookup.scala 33:37]
  assign _T_382 = _T_100 ? 3'h0 : _T_381; // @[Lookup.scala 33:37]
  assign _T_383 = _T_98 ? 3'h0 : _T_382; // @[Lookup.scala 33:37]
  assign _T_384 = _T_96 ? 3'h0 : _T_383; // @[Lookup.scala 33:37]
  assign _T_385 = _T_94 ? 3'h0 : _T_384; // @[Lookup.scala 33:37]
  assign _T_386 = _T_92 ? 3'h0 : _T_385; // @[Lookup.scala 33:37]
  assign _T_387 = _T_90 ? 3'h0 : _T_386; // @[Lookup.scala 33:37]
  assign _T_388 = _T_88 ? 3'h0 : _T_387; // @[Lookup.scala 33:37]
  assign _T_389 = _T_86 ? 3'h0 : _T_388; // @[Lookup.scala 33:37]
  assign _T_390 = _T_84 ? 3'h0 : _T_389; // @[Lookup.scala 33:37]
  assign _T_391 = _T_82 ? 3'h0 : _T_390; // @[Lookup.scala 33:37]
  assign _T_392 = _T_80 ? 3'h0 : _T_391; // @[Lookup.scala 33:37]
  assign _T_393 = _T_78 ? 3'h0 : _T_392; // @[Lookup.scala 33:37]
  assign _T_394 = _T_76 ? 3'h0 : _T_393; // @[Lookup.scala 33:37]
  assign _T_395 = _T_74 ? 3'h0 : _T_394; // @[Lookup.scala 33:37]
  assign _T_396 = _T_72 ? 3'h0 : _T_395; // @[Lookup.scala 33:37]
  assign _T_397 = _T_70 ? 3'h0 : _T_396; // @[Lookup.scala 33:37]
  assign _T_398 = _T_68 ? 3'h0 : _T_397; // @[Lookup.scala 33:37]
  assign _T_399 = _T_66 ? 3'h1 : _T_398; // @[Lookup.scala 33:37]
  assign _T_400 = _T_64 ? 3'h1 : _T_399; // @[Lookup.scala 33:37]
  assign _T_401 = _T_62 ? 3'h1 : _T_400; // @[Lookup.scala 33:37]
  assign _T_402 = _T_60 ? 3'h1 : _T_401; // @[Lookup.scala 33:37]
  assign csignals_5 = _T_58 ? 3'h1 : _T_402; // @[Lookup.scala 33:37]
  assign _T_439 = _T_72 ? 3'h1 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_440 = _T_70 ? 3'h2 : _T_439; // @[Lookup.scala 33:37]
  assign _T_441 = _T_68 ? 3'h3 : _T_440; // @[Lookup.scala 33:37]
  assign _T_442 = _T_66 ? 3'h4 : _T_441; // @[Lookup.scala 33:37]
  assign _T_443 = _T_64 ? 3'h5 : _T_442; // @[Lookup.scala 33:37]
  assign _T_444 = _T_62 ? 3'h1 : _T_443; // @[Lookup.scala 33:37]
  assign _T_445 = _T_60 ? 3'h2 : _T_444; // @[Lookup.scala 33:37]
  assign _T_561 = op2_data == 32'h22; // @[Core.scala 166:55]
  assign _T_562 = _T_557 & _T_561; // @[Core.scala 166:43]
  assign _T_564 = csignals_5 == 3'h1; // @[Core.scala 176:17]
  assign _T_565 = csignals_5 == 3'h2; // @[Core.scala 177:17]
  assign _T_566 = _T_565 ? pc_plus4 : alu_out; // @[Mux.scala 87:16]
  assign io_imem_addr = pc_reg; // @[Core.scala 22:18]
  assign io_dmem_addr = _T_529[31:0]; // @[Core.scala 169:18]
  assign io_dmem_wen = csignals_3[0]; // @[Core.scala 170:17]
  assign io_dmem_wdata = _T_144 ? regfile__T_21_data : _T_27; // @[Core.scala 171:19]
  assign io_dmem_rwtype = _T_58 ? 3'h3 : _T_445; // @[Core.scala 172:20]
  assign io_data = seg_data; // @[Core.scala 165:13]
  initial begin
    $readmemh("/home/star/Desktop/chisel_project/chisel-template/src/main/resources/empty.hex", regfile);
  end
  always @(posedge clock) begin
    if(regfile__T_568_en & regfile__T_568_mask) begin
      regfile[regfile__T_568_addr] <= regfile__T_568_data; // @[Core.scala 17:22]
    end
    if (reset) begin
      pc_reg <= 32'h0;
    end else if (br_flg) begin
      pc_reg <= br_target;
    end else if (_T_5) begin
      pc_reg <= alu_out;
    end else if (!(ecall_flg)) begin
      pc_reg <= pc_plus4;
    end
    if (reset) begin
      seg_data <= 32'h0;
    end else if (_T_562) begin
      if (_T_449) begin
        if (_T_144) begin
          seg_data <= regfile__T_21_data;
        end else if (_T_26) begin
          seg_data <= 32'h0;
        end else begin
          seg_data <= regfile__T_18_data;
        end
      end else if (_T_450) begin
        seg_data <= imm_i_sext;
      end else if (_T_451) begin
        seg_data <= imm_s_sext;
      end else if (_T_452) begin
        seg_data <= imm_j_sext;
      end else if (_T_453) begin
        seg_data <= imm_u_shifted;
      end else begin
        seg_data <= 32'h0;
      end
    end
  end
endmodule
module Rom(
  input         clock,
  input  [31:0] io_addr,
  output [31:0] io_inst
);
  reg [31:0] mem [0:4095]; // @[Rom.scala 17:18]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_2_data; // @[Rom.scala 17:18]
  wire [11:0] mem__T_2_addr; // @[Rom.scala 17:18]
  wire [29:0] _T; // @[Rom.scala 19:27]
  assign mem__T_2_addr = _T[11:0];
  assign mem__T_2_data = mem[mem__T_2_addr]; // @[Rom.scala 17:18]
  assign _T = io_addr[31:2]; // @[Rom.scala 19:27]
  assign io_inst = mem__T_2_data; // @[Rom.scala 19:13]
  initial begin
    $readmemh("/home/star/Desktop/chisel_project/chisel-template/src/main/resources/risc-v-benchmark_ccab.hex", mem);
  end
endmodule
module Ram(
  input         clock,
  input  [31:0] io_addr,
  output [31:0] io_rdata,
  input         io_wen,
  input  [31:0] io_wdata,
  input  [2:0]  io_rwtype
);
  reg [7:0] mem_0 [0:16383]; // @[Ram.scala 18:18]
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_4_data; // @[Ram.scala 18:18]
  wire [13:0] mem_0__T_4_addr; // @[Ram.scala 18:18]
  wire [7:0] mem_0__T_2_data; // @[Ram.scala 18:18]
  wire [13:0] mem_0__T_2_addr; // @[Ram.scala 18:18]
  wire  mem_0__T_2_mask; // @[Ram.scala 18:18]
  wire  mem_0__T_2_en; // @[Ram.scala 18:18]
  reg [7:0] mem_1 [0:16383]; // @[Ram.scala 18:18]
  reg [31:0] _RAND_1;
  wire [7:0] mem_1__T_4_data; // @[Ram.scala 18:18]
  wire [13:0] mem_1__T_4_addr; // @[Ram.scala 18:18]
  wire [7:0] mem_1__T_2_data; // @[Ram.scala 18:18]
  wire [13:0] mem_1__T_2_addr; // @[Ram.scala 18:18]
  wire  mem_1__T_2_mask; // @[Ram.scala 18:18]
  wire  mem_1__T_2_en; // @[Ram.scala 18:18]
  reg [7:0] mem_2 [0:16383]; // @[Ram.scala 18:18]
  reg [31:0] _RAND_2;
  wire [7:0] mem_2__T_4_data; // @[Ram.scala 18:18]
  wire [13:0] mem_2__T_4_addr; // @[Ram.scala 18:18]
  wire [7:0] mem_2__T_2_data; // @[Ram.scala 18:18]
  wire [13:0] mem_2__T_2_addr; // @[Ram.scala 18:18]
  wire  mem_2__T_2_mask; // @[Ram.scala 18:18]
  wire  mem_2__T_2_en; // @[Ram.scala 18:18]
  reg [7:0] mem_3 [0:16383]; // @[Ram.scala 18:18]
  reg [31:0] _RAND_3;
  wire [7:0] mem_3__T_4_data; // @[Ram.scala 18:18]
  wire [13:0] mem_3__T_4_addr; // @[Ram.scala 18:18]
  wire [7:0] mem_3__T_2_data; // @[Ram.scala 18:18]
  wire [13:0] mem_3__T_2_addr; // @[Ram.scala 18:18]
  wire  mem_3__T_2_mask; // @[Ram.scala 18:18]
  wire  mem_3__T_2_en; // @[Ram.scala 18:18]
  wire [29:0] _T; // @[Ram.scala 25:26]
  wire  _T_5; // @[Ram.scala 34:24]
  wire  _T_7; // @[Ram.scala 38:28]
  wire  _T_8; // @[Ram.scala 38:50]
  wire  _T_9; // @[Ram.scala 38:37]
  wire [1:0] _T_11; // @[Ram.scala 40:36]
  wire  _T_12; // @[Ram.scala 40:53]
  wire  _T_13; // @[Ram.scala 42:32]
  wire  _T_14; // @[Ram.scala 42:54]
  wire  _T_15; // @[Ram.scala 42:41]
  wire  _T_17; // @[Ram.scala 44:39]
  wire  _GEN_25; // @[Ram.scala 42:65]
  wire  _GEN_27; // @[Ram.scala 38:61]
  wire [7:0] _T_6; // @[Ram.scala 35:39]
  wire [7:0] _GEN_24; // @[Ram.scala 42:65]
  wire [7:0] _GEN_26; // @[Ram.scala 38:61]
  wire  _T_26; // @[Ram.scala 40:53]
  wire  _GEN_33; // @[Ram.scala 38:61]
  wire [7:0] _T_20; // @[Ram.scala 35:39]
  wire [7:0] _GEN_30; // @[Ram.scala 42:65]
  wire [7:0] _GEN_32; // @[Ram.scala 38:61]
  wire  _T_40; // @[Ram.scala 40:53]
  wire  _GEN_39; // @[Ram.scala 38:61]
  wire [7:0] _T_34; // @[Ram.scala 35:39]
  wire  _T_54; // @[Ram.scala 40:53]
  wire  _GEN_45; // @[Ram.scala 38:61]
  wire [7:0] _T_48; // @[Ram.scala 35:39]
  wire [7:0] dataOut_temp_0; // @[Ram.scala 24:19]
  wire [7:0] dataOut_temp_1; // @[Ram.scala 24:19]
  wire [7:0] dataOut_temp_2; // @[Ram.scala 24:19]
  wire [7:0] dataOut_temp_3; // @[Ram.scala 24:19]
  wire [31:0] _T_64; // @[Cat.scala 29:58]
  wire [7:0] _GEN_49; // @[Ram.scala 55:73]
  wire [7:0] _GEN_50; // @[Ram.scala 55:73]
  wire [7:0] _GEN_51; // @[Ram.scala 55:73]
  wire  _T_67; // @[Ram.scala 55:73]
  wire [23:0] _T_69; // @[Bitwise.scala 71:12]
  wire [31:0] _T_71; // @[Cat.scala 29:58]
  wire [103:0] _T_74; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[Ram.scala 57:72]
  wire [7:0] _GEN_61; // @[Ram.scala 57:78]
  wire [7:0] _GEN_62; // @[Ram.scala 57:78]
  wire [7:0] _GEN_63; // @[Ram.scala 57:78]
  wire  _T_79; // @[Ram.scala 57:78]
  wire [15:0] _T_81; // @[Bitwise.scala 71:12]
  wire [31:0] _T_87; // @[Cat.scala 29:58]
  wire [79:0] _T_94; // @[Cat.scala 29:58]
  wire [79:0] _T_95; // @[Mux.scala 87:16]
  wire [79:0] _T_96; // @[Mux.scala 87:16]
  wire [103:0] _T_97; // @[Mux.scala 87:16]
  wire [103:0] _T_98; // @[Mux.scala 87:16]
  wire [103:0] _T_99; // @[Mux.scala 87:16]
  assign mem_0__T_4_addr = io_addr[13:0];
  assign mem_0__T_4_data = mem_0[mem_0__T_4_addr]; // @[Ram.scala 18:18]
  assign mem_0__T_2_data = _T_5 ? _T_6 : _GEN_26;
  assign mem_0__T_2_addr = _T[13:0];
  assign mem_0__T_2_mask = _T_5 | _GEN_27;
  assign mem_0__T_2_en = io_wen;
  assign mem_1__T_4_addr = io_addr[13:0];
  assign mem_1__T_4_data = mem_1[mem_1__T_4_addr]; // @[Ram.scala 18:18]
  assign mem_1__T_2_data = _T_5 ? _T_20 : _GEN_32;
  assign mem_1__T_2_addr = _T[13:0];
  assign mem_1__T_2_mask = _T_5 | _GEN_33;
  assign mem_1__T_2_en = io_wen;
  assign mem_2__T_4_addr = io_addr[13:0];
  assign mem_2__T_4_data = mem_2[mem_2__T_4_addr]; // @[Ram.scala 18:18]
  assign mem_2__T_2_data = _T_5 ? _T_34 : _GEN_26;
  assign mem_2__T_2_addr = _T[13:0];
  assign mem_2__T_2_mask = _T_5 | _GEN_39;
  assign mem_2__T_2_en = io_wen;
  assign mem_3__T_4_addr = io_addr[13:0];
  assign mem_3__T_4_data = mem_3[mem_3__T_4_addr]; // @[Ram.scala 18:18]
  assign mem_3__T_2_data = _T_5 ? _T_48 : _GEN_32;
  assign mem_3__T_2_addr = _T[13:0];
  assign mem_3__T_2_mask = _T_5 | _GEN_45;
  assign mem_3__T_2_en = io_wen;
  assign _T = io_addr[31:2]; // @[Ram.scala 25:26]
  assign _T_5 = io_rwtype == 3'h1; // @[Ram.scala 34:24]
  assign _T_7 = io_rwtype == 3'h3; // @[Ram.scala 38:28]
  assign _T_8 = io_rwtype == 3'h5; // @[Ram.scala 38:50]
  assign _T_9 = _T_7 | _T_8; // @[Ram.scala 38:37]
  assign _T_11 = io_addr[1:0]; // @[Ram.scala 40:36]
  assign _T_12 = _T_11 == 2'h0; // @[Ram.scala 40:53]
  assign _T_13 = io_rwtype == 3'h2; // @[Ram.scala 42:32]
  assign _T_14 = io_rwtype == 3'h4; // @[Ram.scala 42:54]
  assign _T_15 = _T_13 | _T_14; // @[Ram.scala 42:41]
  assign _T_17 = io_addr[1]; // @[Ram.scala 44:39]
  assign _GEN_25 = _T_15 & _T_17; // @[Ram.scala 42:65]
  assign _GEN_27 = _T_9 ? _T_12 : _GEN_25; // @[Ram.scala 38:61]
  assign _T_6 = io_wdata[7:0]; // @[Ram.scala 35:39]
  assign _GEN_24 = _T_15 ? _T_6 : 8'h0; // @[Ram.scala 42:65]
  assign _GEN_26 = _T_9 ? _T_6 : _GEN_24; // @[Ram.scala 38:61]
  assign _T_26 = _T_11 == 2'h1; // @[Ram.scala 40:53]
  assign _GEN_33 = _T_9 ? _T_26 : _GEN_25; // @[Ram.scala 38:61]
  assign _T_20 = io_wdata[15:8]; // @[Ram.scala 35:39]
  assign _GEN_30 = _T_15 ? _T_20 : 8'h0; // @[Ram.scala 42:65]
  assign _GEN_32 = _T_9 ? _T_6 : _GEN_30; // @[Ram.scala 38:61]
  assign _T_40 = _T_11 == 2'h2; // @[Ram.scala 40:53]
  assign _GEN_39 = _T_9 ? _T_40 : _GEN_25; // @[Ram.scala 38:61]
  assign _T_34 = io_wdata[23:16]; // @[Ram.scala 35:39]
  assign _T_54 = _T_11 == 2'h3; // @[Ram.scala 40:53]
  assign _GEN_45 = _T_9 ? _T_54 : _GEN_25; // @[Ram.scala 38:61]
  assign _T_48 = io_wdata[31:24]; // @[Ram.scala 35:39]
  assign dataOut_temp_0 = io_wen ? mem_0__T_4_data : 8'h0; // @[Ram.scala 24:19]
  assign dataOut_temp_1 = io_wen ? mem_1__T_4_data : 8'h0; // @[Ram.scala 24:19]
  assign dataOut_temp_2 = io_wen ? mem_2__T_4_data : 8'h0; // @[Ram.scala 24:19]
  assign dataOut_temp_3 = io_wen ? mem_3__T_4_data : 8'h0; // @[Ram.scala 24:19]
  assign _T_64 = {dataOut_temp_3,dataOut_temp_2,dataOut_temp_1,dataOut_temp_0}; // @[Cat.scala 29:58]
  assign _GEN_49 = 2'h1 == _T_11 ? dataOut_temp_1 : dataOut_temp_0; // @[Ram.scala 55:73]
  assign _GEN_50 = 2'h2 == _T_11 ? dataOut_temp_2 : _GEN_49; // @[Ram.scala 55:73]
  assign _GEN_51 = 2'h3 == _T_11 ? dataOut_temp_3 : _GEN_50; // @[Ram.scala 55:73]
  assign _T_67 = _GEN_51[7]; // @[Ram.scala 55:73]
  assign _T_69 = _T_67 ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_71 = {_T_69,_GEN_51}; // @[Cat.scala 29:58]
  assign _T_74 = {96'h0,_GEN_51}; // @[Cat.scala 29:58]
  assign _T_78 = _T_11 + 2'h1; // @[Ram.scala 57:72]
  assign _GEN_61 = 2'h1 == _T_78 ? dataOut_temp_1 : dataOut_temp_0; // @[Ram.scala 57:78]
  assign _GEN_62 = 2'h2 == _T_78 ? dataOut_temp_2 : _GEN_61; // @[Ram.scala 57:78]
  assign _GEN_63 = 2'h3 == _T_78 ? dataOut_temp_3 : _GEN_62; // @[Ram.scala 57:78]
  assign _T_79 = _GEN_63[7]; // @[Ram.scala 57:78]
  assign _T_81 = _T_79 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_87 = {_T_81,_GEN_63,_GEN_51}; // @[Cat.scala 29:58]
  assign _T_94 = {64'h0,_GEN_63,_GEN_51}; // @[Cat.scala 29:58]
  assign _T_95 = _T_14 ? _T_94 : 80'h0; // @[Mux.scala 87:16]
  assign _T_96 = _T_13 ? {{48'd0}, _T_87} : _T_95; // @[Mux.scala 87:16]
  assign _T_97 = _T_8 ? _T_74 : {{24'd0}, _T_96}; // @[Mux.scala 87:16]
  assign _T_98 = _T_7 ? {{72'd0}, _T_71} : _T_97; // @[Mux.scala 87:16]
  assign _T_99 = _T_5 ? {{72'd0}, _T_64} : _T_98; // @[Mux.scala 87:16]
  assign io_rdata = _T_99[31:0]; // @[Ram.scala 53:14]
  initial begin
    $readmemh("/home/star/Desktop/chisel_project/chisel-template/src/main/resources/empty.hex", mem);
  end
  always @(posedge clock) begin
    if(mem_0__T_2_en & mem_0__T_2_mask) begin
      mem_0[mem_0__T_2_addr] <= mem_0__T_2_data; // @[Ram.scala 18:18]
    end
    if(mem_1__T_2_en & mem_1__T_2_mask) begin
      mem_1[mem_1__T_2_addr] <= mem_1__T_2_data; // @[Ram.scala 18:18]
    end
    if(mem_2__T_2_en & mem_2__T_2_mask) begin
      mem_2[mem_2__T_2_addr] <= mem_2__T_2_data; // @[Ram.scala 18:18]
    end
    if(mem_3__T_2_en & mem_3__T_2_mask) begin
      mem_3[mem_3__T_2_addr] <= mem_3__T_2_data; // @[Ram.scala 18:18]
    end
  end
endmodule
module Seg(
  input  [31:0] io_data,
  output [7:0]  io_led_0,
  output [7:0]  io_led_1,
  output [7:0]  io_led_2,
  output [7:0]  io_led_3,
  output [7:0]  io_led_4,
  output [7:0]  io_led_5,
  output [7:0]  io_led_6,
  output [7:0]  io_led_7
);
  wire [3:0] _T; // @[Seg.scala 16:21]
  wire  _T_1; // @[Seg.scala 16:40]
  wire  _T_3; // @[Seg.scala 17:40]
  wire  _T_5; // @[Seg.scala 18:40]
  wire  _T_7; // @[Seg.scala 19:40]
  wire  _T_9; // @[Seg.scala 20:40]
  wire  _T_11; // @[Seg.scala 21:40]
  wire  _T_13; // @[Seg.scala 22:40]
  wire  _T_15; // @[Seg.scala 23:40]
  wire  _T_17; // @[Seg.scala 24:40]
  wire  _T_19; // @[Seg.scala 25:40]
  wire  _T_21; // @[Seg.scala 26:40]
  wire  _T_23; // @[Seg.scala 27:40]
  wire  _T_25; // @[Seg.scala 28:40]
  wire  _T_27; // @[Seg.scala 29:40]
  wire  _T_29; // @[Seg.scala 30:40]
  wire [7:0] _T_30; // @[Mux.scala 87:16]
  wire [7:0] _T_31; // @[Mux.scala 87:16]
  wire [7:0] _T_32; // @[Mux.scala 87:16]
  wire [7:0] _T_33; // @[Mux.scala 87:16]
  wire [7:0] _T_34; // @[Mux.scala 87:16]
  wire [7:0] _T_35; // @[Mux.scala 87:16]
  wire [7:0] _T_36; // @[Mux.scala 87:16]
  wire [7:0] _T_37; // @[Mux.scala 87:16]
  wire [7:0] _T_38; // @[Mux.scala 87:16]
  wire [7:0] _T_39; // @[Mux.scala 87:16]
  wire [7:0] _T_40; // @[Mux.scala 87:16]
  wire [7:0] _T_41; // @[Mux.scala 87:16]
  wire [7:0] _T_42; // @[Mux.scala 87:16]
  wire [7:0] _T_43; // @[Mux.scala 87:16]
  wire [3:0] _T_45; // @[Seg.scala 16:21]
  wire  _T_46; // @[Seg.scala 16:40]
  wire  _T_48; // @[Seg.scala 17:40]
  wire  _T_50; // @[Seg.scala 18:40]
  wire  _T_52; // @[Seg.scala 19:40]
  wire  _T_54; // @[Seg.scala 20:40]
  wire  _T_56; // @[Seg.scala 21:40]
  wire  _T_58; // @[Seg.scala 22:40]
  wire  _T_60; // @[Seg.scala 23:40]
  wire  _T_62; // @[Seg.scala 24:40]
  wire  _T_64; // @[Seg.scala 25:40]
  wire  _T_66; // @[Seg.scala 26:40]
  wire  _T_68; // @[Seg.scala 27:40]
  wire  _T_70; // @[Seg.scala 28:40]
  wire  _T_72; // @[Seg.scala 29:40]
  wire  _T_74; // @[Seg.scala 30:40]
  wire [7:0] _T_75; // @[Mux.scala 87:16]
  wire [7:0] _T_76; // @[Mux.scala 87:16]
  wire [7:0] _T_77; // @[Mux.scala 87:16]
  wire [7:0] _T_78; // @[Mux.scala 87:16]
  wire [7:0] _T_79; // @[Mux.scala 87:16]
  wire [7:0] _T_80; // @[Mux.scala 87:16]
  wire [7:0] _T_81; // @[Mux.scala 87:16]
  wire [7:0] _T_82; // @[Mux.scala 87:16]
  wire [7:0] _T_83; // @[Mux.scala 87:16]
  wire [7:0] _T_84; // @[Mux.scala 87:16]
  wire [7:0] _T_85; // @[Mux.scala 87:16]
  wire [7:0] _T_86; // @[Mux.scala 87:16]
  wire [7:0] _T_87; // @[Mux.scala 87:16]
  wire [7:0] _T_88; // @[Mux.scala 87:16]
  wire [3:0] _T_90; // @[Seg.scala 16:21]
  wire  _T_91; // @[Seg.scala 16:40]
  wire  _T_93; // @[Seg.scala 17:40]
  wire  _T_95; // @[Seg.scala 18:40]
  wire  _T_97; // @[Seg.scala 19:40]
  wire  _T_99; // @[Seg.scala 20:40]
  wire  _T_101; // @[Seg.scala 21:40]
  wire  _T_103; // @[Seg.scala 22:40]
  wire  _T_105; // @[Seg.scala 23:40]
  wire  _T_107; // @[Seg.scala 24:40]
  wire  _T_109; // @[Seg.scala 25:40]
  wire  _T_111; // @[Seg.scala 26:40]
  wire  _T_113; // @[Seg.scala 27:40]
  wire  _T_115; // @[Seg.scala 28:40]
  wire  _T_117; // @[Seg.scala 29:40]
  wire  _T_119; // @[Seg.scala 30:40]
  wire [7:0] _T_120; // @[Mux.scala 87:16]
  wire [7:0] _T_121; // @[Mux.scala 87:16]
  wire [7:0] _T_122; // @[Mux.scala 87:16]
  wire [7:0] _T_123; // @[Mux.scala 87:16]
  wire [7:0] _T_124; // @[Mux.scala 87:16]
  wire [7:0] _T_125; // @[Mux.scala 87:16]
  wire [7:0] _T_126; // @[Mux.scala 87:16]
  wire [7:0] _T_127; // @[Mux.scala 87:16]
  wire [7:0] _T_128; // @[Mux.scala 87:16]
  wire [7:0] _T_129; // @[Mux.scala 87:16]
  wire [7:0] _T_130; // @[Mux.scala 87:16]
  wire [7:0] _T_131; // @[Mux.scala 87:16]
  wire [7:0] _T_132; // @[Mux.scala 87:16]
  wire [7:0] _T_133; // @[Mux.scala 87:16]
  wire [3:0] _T_135; // @[Seg.scala 16:21]
  wire  _T_136; // @[Seg.scala 16:40]
  wire  _T_138; // @[Seg.scala 17:40]
  wire  _T_140; // @[Seg.scala 18:40]
  wire  _T_142; // @[Seg.scala 19:40]
  wire  _T_144; // @[Seg.scala 20:40]
  wire  _T_146; // @[Seg.scala 21:40]
  wire  _T_148; // @[Seg.scala 22:40]
  wire  _T_150; // @[Seg.scala 23:40]
  wire  _T_152; // @[Seg.scala 24:40]
  wire  _T_154; // @[Seg.scala 25:40]
  wire  _T_156; // @[Seg.scala 26:40]
  wire  _T_158; // @[Seg.scala 27:40]
  wire  _T_160; // @[Seg.scala 28:40]
  wire  _T_162; // @[Seg.scala 29:40]
  wire  _T_164; // @[Seg.scala 30:40]
  wire [7:0] _T_165; // @[Mux.scala 87:16]
  wire [7:0] _T_166; // @[Mux.scala 87:16]
  wire [7:0] _T_167; // @[Mux.scala 87:16]
  wire [7:0] _T_168; // @[Mux.scala 87:16]
  wire [7:0] _T_169; // @[Mux.scala 87:16]
  wire [7:0] _T_170; // @[Mux.scala 87:16]
  wire [7:0] _T_171; // @[Mux.scala 87:16]
  wire [7:0] _T_172; // @[Mux.scala 87:16]
  wire [7:0] _T_173; // @[Mux.scala 87:16]
  wire [7:0] _T_174; // @[Mux.scala 87:16]
  wire [7:0] _T_175; // @[Mux.scala 87:16]
  wire [7:0] _T_176; // @[Mux.scala 87:16]
  wire [7:0] _T_177; // @[Mux.scala 87:16]
  wire [7:0] _T_178; // @[Mux.scala 87:16]
  wire [3:0] _T_180; // @[Seg.scala 16:21]
  wire  _T_181; // @[Seg.scala 16:40]
  wire  _T_183; // @[Seg.scala 17:40]
  wire  _T_185; // @[Seg.scala 18:40]
  wire  _T_187; // @[Seg.scala 19:40]
  wire  _T_189; // @[Seg.scala 20:40]
  wire  _T_191; // @[Seg.scala 21:40]
  wire  _T_193; // @[Seg.scala 22:40]
  wire  _T_195; // @[Seg.scala 23:40]
  wire  _T_197; // @[Seg.scala 24:40]
  wire  _T_199; // @[Seg.scala 25:40]
  wire  _T_201; // @[Seg.scala 26:40]
  wire  _T_203; // @[Seg.scala 27:40]
  wire  _T_205; // @[Seg.scala 28:40]
  wire  _T_207; // @[Seg.scala 29:40]
  wire  _T_209; // @[Seg.scala 30:40]
  wire [7:0] _T_210; // @[Mux.scala 87:16]
  wire [7:0] _T_211; // @[Mux.scala 87:16]
  wire [7:0] _T_212; // @[Mux.scala 87:16]
  wire [7:0] _T_213; // @[Mux.scala 87:16]
  wire [7:0] _T_214; // @[Mux.scala 87:16]
  wire [7:0] _T_215; // @[Mux.scala 87:16]
  wire [7:0] _T_216; // @[Mux.scala 87:16]
  wire [7:0] _T_217; // @[Mux.scala 87:16]
  wire [7:0] _T_218; // @[Mux.scala 87:16]
  wire [7:0] _T_219; // @[Mux.scala 87:16]
  wire [7:0] _T_220; // @[Mux.scala 87:16]
  wire [7:0] _T_221; // @[Mux.scala 87:16]
  wire [7:0] _T_222; // @[Mux.scala 87:16]
  wire [7:0] _T_223; // @[Mux.scala 87:16]
  wire [3:0] _T_225; // @[Seg.scala 16:21]
  wire  _T_226; // @[Seg.scala 16:40]
  wire  _T_228; // @[Seg.scala 17:40]
  wire  _T_230; // @[Seg.scala 18:40]
  wire  _T_232; // @[Seg.scala 19:40]
  wire  _T_234; // @[Seg.scala 20:40]
  wire  _T_236; // @[Seg.scala 21:40]
  wire  _T_238; // @[Seg.scala 22:40]
  wire  _T_240; // @[Seg.scala 23:40]
  wire  _T_242; // @[Seg.scala 24:40]
  wire  _T_244; // @[Seg.scala 25:40]
  wire  _T_246; // @[Seg.scala 26:40]
  wire  _T_248; // @[Seg.scala 27:40]
  wire  _T_250; // @[Seg.scala 28:40]
  wire  _T_252; // @[Seg.scala 29:40]
  wire  _T_254; // @[Seg.scala 30:40]
  wire [7:0] _T_255; // @[Mux.scala 87:16]
  wire [7:0] _T_256; // @[Mux.scala 87:16]
  wire [7:0] _T_257; // @[Mux.scala 87:16]
  wire [7:0] _T_258; // @[Mux.scala 87:16]
  wire [7:0] _T_259; // @[Mux.scala 87:16]
  wire [7:0] _T_260; // @[Mux.scala 87:16]
  wire [7:0] _T_261; // @[Mux.scala 87:16]
  wire [7:0] _T_262; // @[Mux.scala 87:16]
  wire [7:0] _T_263; // @[Mux.scala 87:16]
  wire [7:0] _T_264; // @[Mux.scala 87:16]
  wire [7:0] _T_265; // @[Mux.scala 87:16]
  wire [7:0] _T_266; // @[Mux.scala 87:16]
  wire [7:0] _T_267; // @[Mux.scala 87:16]
  wire [7:0] _T_268; // @[Mux.scala 87:16]
  wire [3:0] _T_270; // @[Seg.scala 16:21]
  wire  _T_271; // @[Seg.scala 16:40]
  wire  _T_273; // @[Seg.scala 17:40]
  wire  _T_275; // @[Seg.scala 18:40]
  wire  _T_277; // @[Seg.scala 19:40]
  wire  _T_279; // @[Seg.scala 20:40]
  wire  _T_281; // @[Seg.scala 21:40]
  wire  _T_283; // @[Seg.scala 22:40]
  wire  _T_285; // @[Seg.scala 23:40]
  wire  _T_287; // @[Seg.scala 24:40]
  wire  _T_289; // @[Seg.scala 25:40]
  wire  _T_291; // @[Seg.scala 26:40]
  wire  _T_293; // @[Seg.scala 27:40]
  wire  _T_295; // @[Seg.scala 28:40]
  wire  _T_297; // @[Seg.scala 29:40]
  wire  _T_299; // @[Seg.scala 30:40]
  wire [7:0] _T_300; // @[Mux.scala 87:16]
  wire [7:0] _T_301; // @[Mux.scala 87:16]
  wire [7:0] _T_302; // @[Mux.scala 87:16]
  wire [7:0] _T_303; // @[Mux.scala 87:16]
  wire [7:0] _T_304; // @[Mux.scala 87:16]
  wire [7:0] _T_305; // @[Mux.scala 87:16]
  wire [7:0] _T_306; // @[Mux.scala 87:16]
  wire [7:0] _T_307; // @[Mux.scala 87:16]
  wire [7:0] _T_308; // @[Mux.scala 87:16]
  wire [7:0] _T_309; // @[Mux.scala 87:16]
  wire [7:0] _T_310; // @[Mux.scala 87:16]
  wire [7:0] _T_311; // @[Mux.scala 87:16]
  wire [7:0] _T_312; // @[Mux.scala 87:16]
  wire [7:0] _T_313; // @[Mux.scala 87:16]
  wire [3:0] _T_315; // @[Seg.scala 16:21]
  wire  _T_316; // @[Seg.scala 16:40]
  wire  _T_318; // @[Seg.scala 17:40]
  wire  _T_320; // @[Seg.scala 18:40]
  wire  _T_322; // @[Seg.scala 19:40]
  wire  _T_324; // @[Seg.scala 20:40]
  wire  _T_326; // @[Seg.scala 21:40]
  wire  _T_328; // @[Seg.scala 22:40]
  wire  _T_330; // @[Seg.scala 23:40]
  wire  _T_332; // @[Seg.scala 24:40]
  wire  _T_334; // @[Seg.scala 25:40]
  wire  _T_336; // @[Seg.scala 26:40]
  wire  _T_338; // @[Seg.scala 27:40]
  wire  _T_340; // @[Seg.scala 28:40]
  wire  _T_342; // @[Seg.scala 29:40]
  wire  _T_344; // @[Seg.scala 30:40]
  wire [7:0] _T_345; // @[Mux.scala 87:16]
  wire [7:0] _T_346; // @[Mux.scala 87:16]
  wire [7:0] _T_347; // @[Mux.scala 87:16]
  wire [7:0] _T_348; // @[Mux.scala 87:16]
  wire [7:0] _T_349; // @[Mux.scala 87:16]
  wire [7:0] _T_350; // @[Mux.scala 87:16]
  wire [7:0] _T_351; // @[Mux.scala 87:16]
  wire [7:0] _T_352; // @[Mux.scala 87:16]
  wire [7:0] _T_353; // @[Mux.scala 87:16]
  wire [7:0] _T_354; // @[Mux.scala 87:16]
  wire [7:0] _T_355; // @[Mux.scala 87:16]
  wire [7:0] _T_356; // @[Mux.scala 87:16]
  wire [7:0] _T_357; // @[Mux.scala 87:16]
  wire [7:0] _T_358; // @[Mux.scala 87:16]
  assign _T = io_data[3:0]; // @[Seg.scala 16:21]
  assign _T_1 = _T == 4'h0; // @[Seg.scala 16:40]
  assign _T_3 = _T == 4'h1; // @[Seg.scala 17:40]
  assign _T_5 = _T == 4'h2; // @[Seg.scala 18:40]
  assign _T_7 = _T == 4'h3; // @[Seg.scala 19:40]
  assign _T_9 = _T == 4'h4; // @[Seg.scala 20:40]
  assign _T_11 = _T == 4'h5; // @[Seg.scala 21:40]
  assign _T_13 = _T == 4'h6; // @[Seg.scala 22:40]
  assign _T_15 = _T == 4'h7; // @[Seg.scala 23:40]
  assign _T_17 = _T == 4'h8; // @[Seg.scala 24:40]
  assign _T_19 = _T == 4'h9; // @[Seg.scala 25:40]
  assign _T_21 = _T == 4'ha; // @[Seg.scala 26:40]
  assign _T_23 = _T == 4'hb; // @[Seg.scala 27:40]
  assign _T_25 = _T == 4'hc; // @[Seg.scala 28:40]
  assign _T_27 = _T == 4'hd; // @[Seg.scala 29:40]
  assign _T_29 = _T == 4'he; // @[Seg.scala 30:40]
  assign _T_30 = _T_29 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_31 = _T_27 ? 8'ha1 : _T_30; // @[Mux.scala 87:16]
  assign _T_32 = _T_25 ? 8'hc6 : _T_31; // @[Mux.scala 87:16]
  assign _T_33 = _T_23 ? 8'h83 : _T_32; // @[Mux.scala 87:16]
  assign _T_34 = _T_21 ? 8'h88 : _T_33; // @[Mux.scala 87:16]
  assign _T_35 = _T_19 ? 8'h98 : _T_34; // @[Mux.scala 87:16]
  assign _T_36 = _T_17 ? 8'h80 : _T_35; // @[Mux.scala 87:16]
  assign _T_37 = _T_15 ? 8'hf8 : _T_36; // @[Mux.scala 87:16]
  assign _T_38 = _T_13 ? 8'h82 : _T_37; // @[Mux.scala 87:16]
  assign _T_39 = _T_11 ? 8'h92 : _T_38; // @[Mux.scala 87:16]
  assign _T_40 = _T_9 ? 8'h99 : _T_39; // @[Mux.scala 87:16]
  assign _T_41 = _T_7 ? 8'hb0 : _T_40; // @[Mux.scala 87:16]
  assign _T_42 = _T_5 ? 8'ha4 : _T_41; // @[Mux.scala 87:16]
  assign _T_43 = _T_3 ? 8'hf9 : _T_42; // @[Mux.scala 87:16]
  assign _T_45 = io_data[7:4]; // @[Seg.scala 16:21]
  assign _T_46 = _T_45 == 4'h0; // @[Seg.scala 16:40]
  assign _T_48 = _T_45 == 4'h1; // @[Seg.scala 17:40]
  assign _T_50 = _T_45 == 4'h2; // @[Seg.scala 18:40]
  assign _T_52 = _T_45 == 4'h3; // @[Seg.scala 19:40]
  assign _T_54 = _T_45 == 4'h4; // @[Seg.scala 20:40]
  assign _T_56 = _T_45 == 4'h5; // @[Seg.scala 21:40]
  assign _T_58 = _T_45 == 4'h6; // @[Seg.scala 22:40]
  assign _T_60 = _T_45 == 4'h7; // @[Seg.scala 23:40]
  assign _T_62 = _T_45 == 4'h8; // @[Seg.scala 24:40]
  assign _T_64 = _T_45 == 4'h9; // @[Seg.scala 25:40]
  assign _T_66 = _T_45 == 4'ha; // @[Seg.scala 26:40]
  assign _T_68 = _T_45 == 4'hb; // @[Seg.scala 27:40]
  assign _T_70 = _T_45 == 4'hc; // @[Seg.scala 28:40]
  assign _T_72 = _T_45 == 4'hd; // @[Seg.scala 29:40]
  assign _T_74 = _T_45 == 4'he; // @[Seg.scala 30:40]
  assign _T_75 = _T_74 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_76 = _T_72 ? 8'ha1 : _T_75; // @[Mux.scala 87:16]
  assign _T_77 = _T_70 ? 8'hc6 : _T_76; // @[Mux.scala 87:16]
  assign _T_78 = _T_68 ? 8'h83 : _T_77; // @[Mux.scala 87:16]
  assign _T_79 = _T_66 ? 8'h88 : _T_78; // @[Mux.scala 87:16]
  assign _T_80 = _T_64 ? 8'h98 : _T_79; // @[Mux.scala 87:16]
  assign _T_81 = _T_62 ? 8'h80 : _T_80; // @[Mux.scala 87:16]
  assign _T_82 = _T_60 ? 8'hf8 : _T_81; // @[Mux.scala 87:16]
  assign _T_83 = _T_58 ? 8'h82 : _T_82; // @[Mux.scala 87:16]
  assign _T_84 = _T_56 ? 8'h92 : _T_83; // @[Mux.scala 87:16]
  assign _T_85 = _T_54 ? 8'h99 : _T_84; // @[Mux.scala 87:16]
  assign _T_86 = _T_52 ? 8'hb0 : _T_85; // @[Mux.scala 87:16]
  assign _T_87 = _T_50 ? 8'ha4 : _T_86; // @[Mux.scala 87:16]
  assign _T_88 = _T_48 ? 8'hf9 : _T_87; // @[Mux.scala 87:16]
  assign _T_90 = io_data[11:8]; // @[Seg.scala 16:21]
  assign _T_91 = _T_90 == 4'h0; // @[Seg.scala 16:40]
  assign _T_93 = _T_90 == 4'h1; // @[Seg.scala 17:40]
  assign _T_95 = _T_90 == 4'h2; // @[Seg.scala 18:40]
  assign _T_97 = _T_90 == 4'h3; // @[Seg.scala 19:40]
  assign _T_99 = _T_90 == 4'h4; // @[Seg.scala 20:40]
  assign _T_101 = _T_90 == 4'h5; // @[Seg.scala 21:40]
  assign _T_103 = _T_90 == 4'h6; // @[Seg.scala 22:40]
  assign _T_105 = _T_90 == 4'h7; // @[Seg.scala 23:40]
  assign _T_107 = _T_90 == 4'h8; // @[Seg.scala 24:40]
  assign _T_109 = _T_90 == 4'h9; // @[Seg.scala 25:40]
  assign _T_111 = _T_90 == 4'ha; // @[Seg.scala 26:40]
  assign _T_113 = _T_90 == 4'hb; // @[Seg.scala 27:40]
  assign _T_115 = _T_90 == 4'hc; // @[Seg.scala 28:40]
  assign _T_117 = _T_90 == 4'hd; // @[Seg.scala 29:40]
  assign _T_119 = _T_90 == 4'he; // @[Seg.scala 30:40]
  assign _T_120 = _T_119 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_121 = _T_117 ? 8'ha1 : _T_120; // @[Mux.scala 87:16]
  assign _T_122 = _T_115 ? 8'hc6 : _T_121; // @[Mux.scala 87:16]
  assign _T_123 = _T_113 ? 8'h83 : _T_122; // @[Mux.scala 87:16]
  assign _T_124 = _T_111 ? 8'h88 : _T_123; // @[Mux.scala 87:16]
  assign _T_125 = _T_109 ? 8'h98 : _T_124; // @[Mux.scala 87:16]
  assign _T_126 = _T_107 ? 8'h80 : _T_125; // @[Mux.scala 87:16]
  assign _T_127 = _T_105 ? 8'hf8 : _T_126; // @[Mux.scala 87:16]
  assign _T_128 = _T_103 ? 8'h82 : _T_127; // @[Mux.scala 87:16]
  assign _T_129 = _T_101 ? 8'h92 : _T_128; // @[Mux.scala 87:16]
  assign _T_130 = _T_99 ? 8'h99 : _T_129; // @[Mux.scala 87:16]
  assign _T_131 = _T_97 ? 8'hb0 : _T_130; // @[Mux.scala 87:16]
  assign _T_132 = _T_95 ? 8'ha4 : _T_131; // @[Mux.scala 87:16]
  assign _T_133 = _T_93 ? 8'hf9 : _T_132; // @[Mux.scala 87:16]
  assign _T_135 = io_data[15:12]; // @[Seg.scala 16:21]
  assign _T_136 = _T_135 == 4'h0; // @[Seg.scala 16:40]
  assign _T_138 = _T_135 == 4'h1; // @[Seg.scala 17:40]
  assign _T_140 = _T_135 == 4'h2; // @[Seg.scala 18:40]
  assign _T_142 = _T_135 == 4'h3; // @[Seg.scala 19:40]
  assign _T_144 = _T_135 == 4'h4; // @[Seg.scala 20:40]
  assign _T_146 = _T_135 == 4'h5; // @[Seg.scala 21:40]
  assign _T_148 = _T_135 == 4'h6; // @[Seg.scala 22:40]
  assign _T_150 = _T_135 == 4'h7; // @[Seg.scala 23:40]
  assign _T_152 = _T_135 == 4'h8; // @[Seg.scala 24:40]
  assign _T_154 = _T_135 == 4'h9; // @[Seg.scala 25:40]
  assign _T_156 = _T_135 == 4'ha; // @[Seg.scala 26:40]
  assign _T_158 = _T_135 == 4'hb; // @[Seg.scala 27:40]
  assign _T_160 = _T_135 == 4'hc; // @[Seg.scala 28:40]
  assign _T_162 = _T_135 == 4'hd; // @[Seg.scala 29:40]
  assign _T_164 = _T_135 == 4'he; // @[Seg.scala 30:40]
  assign _T_165 = _T_164 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_166 = _T_162 ? 8'ha1 : _T_165; // @[Mux.scala 87:16]
  assign _T_167 = _T_160 ? 8'hc6 : _T_166; // @[Mux.scala 87:16]
  assign _T_168 = _T_158 ? 8'h83 : _T_167; // @[Mux.scala 87:16]
  assign _T_169 = _T_156 ? 8'h88 : _T_168; // @[Mux.scala 87:16]
  assign _T_170 = _T_154 ? 8'h98 : _T_169; // @[Mux.scala 87:16]
  assign _T_171 = _T_152 ? 8'h80 : _T_170; // @[Mux.scala 87:16]
  assign _T_172 = _T_150 ? 8'hf8 : _T_171; // @[Mux.scala 87:16]
  assign _T_173 = _T_148 ? 8'h82 : _T_172; // @[Mux.scala 87:16]
  assign _T_174 = _T_146 ? 8'h92 : _T_173; // @[Mux.scala 87:16]
  assign _T_175 = _T_144 ? 8'h99 : _T_174; // @[Mux.scala 87:16]
  assign _T_176 = _T_142 ? 8'hb0 : _T_175; // @[Mux.scala 87:16]
  assign _T_177 = _T_140 ? 8'ha4 : _T_176; // @[Mux.scala 87:16]
  assign _T_178 = _T_138 ? 8'hf9 : _T_177; // @[Mux.scala 87:16]
  assign _T_180 = io_data[19:16]; // @[Seg.scala 16:21]
  assign _T_181 = _T_180 == 4'h0; // @[Seg.scala 16:40]
  assign _T_183 = _T_180 == 4'h1; // @[Seg.scala 17:40]
  assign _T_185 = _T_180 == 4'h2; // @[Seg.scala 18:40]
  assign _T_187 = _T_180 == 4'h3; // @[Seg.scala 19:40]
  assign _T_189 = _T_180 == 4'h4; // @[Seg.scala 20:40]
  assign _T_191 = _T_180 == 4'h5; // @[Seg.scala 21:40]
  assign _T_193 = _T_180 == 4'h6; // @[Seg.scala 22:40]
  assign _T_195 = _T_180 == 4'h7; // @[Seg.scala 23:40]
  assign _T_197 = _T_180 == 4'h8; // @[Seg.scala 24:40]
  assign _T_199 = _T_180 == 4'h9; // @[Seg.scala 25:40]
  assign _T_201 = _T_180 == 4'ha; // @[Seg.scala 26:40]
  assign _T_203 = _T_180 == 4'hb; // @[Seg.scala 27:40]
  assign _T_205 = _T_180 == 4'hc; // @[Seg.scala 28:40]
  assign _T_207 = _T_180 == 4'hd; // @[Seg.scala 29:40]
  assign _T_209 = _T_180 == 4'he; // @[Seg.scala 30:40]
  assign _T_210 = _T_209 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_211 = _T_207 ? 8'ha1 : _T_210; // @[Mux.scala 87:16]
  assign _T_212 = _T_205 ? 8'hc6 : _T_211; // @[Mux.scala 87:16]
  assign _T_213 = _T_203 ? 8'h83 : _T_212; // @[Mux.scala 87:16]
  assign _T_214 = _T_201 ? 8'h88 : _T_213; // @[Mux.scala 87:16]
  assign _T_215 = _T_199 ? 8'h98 : _T_214; // @[Mux.scala 87:16]
  assign _T_216 = _T_197 ? 8'h80 : _T_215; // @[Mux.scala 87:16]
  assign _T_217 = _T_195 ? 8'hf8 : _T_216; // @[Mux.scala 87:16]
  assign _T_218 = _T_193 ? 8'h82 : _T_217; // @[Mux.scala 87:16]
  assign _T_219 = _T_191 ? 8'h92 : _T_218; // @[Mux.scala 87:16]
  assign _T_220 = _T_189 ? 8'h99 : _T_219; // @[Mux.scala 87:16]
  assign _T_221 = _T_187 ? 8'hb0 : _T_220; // @[Mux.scala 87:16]
  assign _T_222 = _T_185 ? 8'ha4 : _T_221; // @[Mux.scala 87:16]
  assign _T_223 = _T_183 ? 8'hf9 : _T_222; // @[Mux.scala 87:16]
  assign _T_225 = io_data[23:20]; // @[Seg.scala 16:21]
  assign _T_226 = _T_225 == 4'h0; // @[Seg.scala 16:40]
  assign _T_228 = _T_225 == 4'h1; // @[Seg.scala 17:40]
  assign _T_230 = _T_225 == 4'h2; // @[Seg.scala 18:40]
  assign _T_232 = _T_225 == 4'h3; // @[Seg.scala 19:40]
  assign _T_234 = _T_225 == 4'h4; // @[Seg.scala 20:40]
  assign _T_236 = _T_225 == 4'h5; // @[Seg.scala 21:40]
  assign _T_238 = _T_225 == 4'h6; // @[Seg.scala 22:40]
  assign _T_240 = _T_225 == 4'h7; // @[Seg.scala 23:40]
  assign _T_242 = _T_225 == 4'h8; // @[Seg.scala 24:40]
  assign _T_244 = _T_225 == 4'h9; // @[Seg.scala 25:40]
  assign _T_246 = _T_225 == 4'ha; // @[Seg.scala 26:40]
  assign _T_248 = _T_225 == 4'hb; // @[Seg.scala 27:40]
  assign _T_250 = _T_225 == 4'hc; // @[Seg.scala 28:40]
  assign _T_252 = _T_225 == 4'hd; // @[Seg.scala 29:40]
  assign _T_254 = _T_225 == 4'he; // @[Seg.scala 30:40]
  assign _T_255 = _T_254 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_256 = _T_252 ? 8'ha1 : _T_255; // @[Mux.scala 87:16]
  assign _T_257 = _T_250 ? 8'hc6 : _T_256; // @[Mux.scala 87:16]
  assign _T_258 = _T_248 ? 8'h83 : _T_257; // @[Mux.scala 87:16]
  assign _T_259 = _T_246 ? 8'h88 : _T_258; // @[Mux.scala 87:16]
  assign _T_260 = _T_244 ? 8'h98 : _T_259; // @[Mux.scala 87:16]
  assign _T_261 = _T_242 ? 8'h80 : _T_260; // @[Mux.scala 87:16]
  assign _T_262 = _T_240 ? 8'hf8 : _T_261; // @[Mux.scala 87:16]
  assign _T_263 = _T_238 ? 8'h82 : _T_262; // @[Mux.scala 87:16]
  assign _T_264 = _T_236 ? 8'h92 : _T_263; // @[Mux.scala 87:16]
  assign _T_265 = _T_234 ? 8'h99 : _T_264; // @[Mux.scala 87:16]
  assign _T_266 = _T_232 ? 8'hb0 : _T_265; // @[Mux.scala 87:16]
  assign _T_267 = _T_230 ? 8'ha4 : _T_266; // @[Mux.scala 87:16]
  assign _T_268 = _T_228 ? 8'hf9 : _T_267; // @[Mux.scala 87:16]
  assign _T_270 = io_data[27:24]; // @[Seg.scala 16:21]
  assign _T_271 = _T_270 == 4'h0; // @[Seg.scala 16:40]
  assign _T_273 = _T_270 == 4'h1; // @[Seg.scala 17:40]
  assign _T_275 = _T_270 == 4'h2; // @[Seg.scala 18:40]
  assign _T_277 = _T_270 == 4'h3; // @[Seg.scala 19:40]
  assign _T_279 = _T_270 == 4'h4; // @[Seg.scala 20:40]
  assign _T_281 = _T_270 == 4'h5; // @[Seg.scala 21:40]
  assign _T_283 = _T_270 == 4'h6; // @[Seg.scala 22:40]
  assign _T_285 = _T_270 == 4'h7; // @[Seg.scala 23:40]
  assign _T_287 = _T_270 == 4'h8; // @[Seg.scala 24:40]
  assign _T_289 = _T_270 == 4'h9; // @[Seg.scala 25:40]
  assign _T_291 = _T_270 == 4'ha; // @[Seg.scala 26:40]
  assign _T_293 = _T_270 == 4'hb; // @[Seg.scala 27:40]
  assign _T_295 = _T_270 == 4'hc; // @[Seg.scala 28:40]
  assign _T_297 = _T_270 == 4'hd; // @[Seg.scala 29:40]
  assign _T_299 = _T_270 == 4'he; // @[Seg.scala 30:40]
  assign _T_300 = _T_299 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_301 = _T_297 ? 8'ha1 : _T_300; // @[Mux.scala 87:16]
  assign _T_302 = _T_295 ? 8'hc6 : _T_301; // @[Mux.scala 87:16]
  assign _T_303 = _T_293 ? 8'h83 : _T_302; // @[Mux.scala 87:16]
  assign _T_304 = _T_291 ? 8'h88 : _T_303; // @[Mux.scala 87:16]
  assign _T_305 = _T_289 ? 8'h98 : _T_304; // @[Mux.scala 87:16]
  assign _T_306 = _T_287 ? 8'h80 : _T_305; // @[Mux.scala 87:16]
  assign _T_307 = _T_285 ? 8'hf8 : _T_306; // @[Mux.scala 87:16]
  assign _T_308 = _T_283 ? 8'h82 : _T_307; // @[Mux.scala 87:16]
  assign _T_309 = _T_281 ? 8'h92 : _T_308; // @[Mux.scala 87:16]
  assign _T_310 = _T_279 ? 8'h99 : _T_309; // @[Mux.scala 87:16]
  assign _T_311 = _T_277 ? 8'hb0 : _T_310; // @[Mux.scala 87:16]
  assign _T_312 = _T_275 ? 8'ha4 : _T_311; // @[Mux.scala 87:16]
  assign _T_313 = _T_273 ? 8'hf9 : _T_312; // @[Mux.scala 87:16]
  assign _T_315 = io_data[31:28]; // @[Seg.scala 16:21]
  assign _T_316 = _T_315 == 4'h0; // @[Seg.scala 16:40]
  assign _T_318 = _T_315 == 4'h1; // @[Seg.scala 17:40]
  assign _T_320 = _T_315 == 4'h2; // @[Seg.scala 18:40]
  assign _T_322 = _T_315 == 4'h3; // @[Seg.scala 19:40]
  assign _T_324 = _T_315 == 4'h4; // @[Seg.scala 20:40]
  assign _T_326 = _T_315 == 4'h5; // @[Seg.scala 21:40]
  assign _T_328 = _T_315 == 4'h6; // @[Seg.scala 22:40]
  assign _T_330 = _T_315 == 4'h7; // @[Seg.scala 23:40]
  assign _T_332 = _T_315 == 4'h8; // @[Seg.scala 24:40]
  assign _T_334 = _T_315 == 4'h9; // @[Seg.scala 25:40]
  assign _T_336 = _T_315 == 4'ha; // @[Seg.scala 26:40]
  assign _T_338 = _T_315 == 4'hb; // @[Seg.scala 27:40]
  assign _T_340 = _T_315 == 4'hc; // @[Seg.scala 28:40]
  assign _T_342 = _T_315 == 4'hd; // @[Seg.scala 29:40]
  assign _T_344 = _T_315 == 4'he; // @[Seg.scala 30:40]
  assign _T_345 = _T_344 ? 8'h86 : 8'h8e; // @[Mux.scala 87:16]
  assign _T_346 = _T_342 ? 8'ha1 : _T_345; // @[Mux.scala 87:16]
  assign _T_347 = _T_340 ? 8'hc6 : _T_346; // @[Mux.scala 87:16]
  assign _T_348 = _T_338 ? 8'h83 : _T_347; // @[Mux.scala 87:16]
  assign _T_349 = _T_336 ? 8'h88 : _T_348; // @[Mux.scala 87:16]
  assign _T_350 = _T_334 ? 8'h98 : _T_349; // @[Mux.scala 87:16]
  assign _T_351 = _T_332 ? 8'h80 : _T_350; // @[Mux.scala 87:16]
  assign _T_352 = _T_330 ? 8'hf8 : _T_351; // @[Mux.scala 87:16]
  assign _T_353 = _T_328 ? 8'h82 : _T_352; // @[Mux.scala 87:16]
  assign _T_354 = _T_326 ? 8'h92 : _T_353; // @[Mux.scala 87:16]
  assign _T_355 = _T_324 ? 8'h99 : _T_354; // @[Mux.scala 87:16]
  assign _T_356 = _T_322 ? 8'hb0 : _T_355; // @[Mux.scala 87:16]
  assign _T_357 = _T_320 ? 8'ha4 : _T_356; // @[Mux.scala 87:16]
  assign _T_358 = _T_318 ? 8'hf9 : _T_357; // @[Mux.scala 87:16]
  assign io_led_0 = _T_1 ? 8'hc0 : _T_43; // @[Seg.scala 15:19]
  assign io_led_1 = _T_46 ? 8'hc0 : _T_88; // @[Seg.scala 15:19]
  assign io_led_2 = _T_91 ? 8'hc0 : _T_133; // @[Seg.scala 15:19]
  assign io_led_3 = _T_136 ? 8'hc0 : _T_178; // @[Seg.scala 15:19]
  assign io_led_4 = _T_181 ? 8'hc0 : _T_223; // @[Seg.scala 15:19]
  assign io_led_5 = _T_226 ? 8'hc0 : _T_268; // @[Seg.scala 15:19]
  assign io_led_6 = _T_271 ? 8'hc0 : _T_313; // @[Seg.scala 15:19]
  assign io_led_7 = _T_316 ? 8'hc0 : _T_358; // @[Seg.scala 15:19]
endmodule
module Top(
  input        clock,
  input        reset,
  output [7:0] io_led_0,
  output [7:0] io_led_1,
  output [7:0] io_led_2,
  output [7:0] io_led_3,
  output [7:0] io_led_4,
  output [7:0] io_led_5,
  output [7:0] io_led_6,
  output [7:0] io_led_7
);
  wire  core_clock; // @[Top.scala 10:22]
  wire  core_reset; // @[Top.scala 10:22]
  wire [31:0] core_io_imem_addr; // @[Top.scala 10:22]
  wire [31:0] core_io_imem_inst; // @[Top.scala 10:22]
  wire [31:0] core_io_dmem_addr; // @[Top.scala 10:22]
  wire [31:0] core_io_dmem_rdata; // @[Top.scala 10:22]
  wire  core_io_dmem_wen; // @[Top.scala 10:22]
  wire [31:0] core_io_dmem_wdata; // @[Top.scala 10:22]
  wire [2:0] core_io_dmem_rwtype; // @[Top.scala 10:22]
  wire [31:0] core_io_data; // @[Top.scala 10:22]
  wire  rom_clock; // @[Top.scala 11:21]
  wire [31:0] rom_io_addr; // @[Top.scala 11:21]
  wire [31:0] rom_io_inst; // @[Top.scala 11:21]
  wire  ram_clock; // @[Top.scala 12:21]
  wire [31:0] ram_io_addr; // @[Top.scala 12:21]
  wire [31:0] ram_io_rdata; // @[Top.scala 12:21]
  wire  ram_io_wen; // @[Top.scala 12:21]
  wire [31:0] ram_io_wdata; // @[Top.scala 12:21]
  wire [2:0] ram_io_rwtype; // @[Top.scala 12:21]
  wire [31:0] seg_io_data; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_0; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_1; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_2; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_3; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_4; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_5; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_6; // @[Top.scala 13:21]
  wire [7:0] seg_io_led_7; // @[Top.scala 13:21]
  Core core ( // @[Top.scala 10:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_addr(core_io_imem_addr),
    .io_imem_inst(core_io_imem_inst),
    .io_dmem_addr(core_io_dmem_addr),
    .io_dmem_rdata(core_io_dmem_rdata),
    .io_dmem_wen(core_io_dmem_wen),
    .io_dmem_wdata(core_io_dmem_wdata),
    .io_dmem_rwtype(core_io_dmem_rwtype),
    .io_data(core_io_data)
  );
  Rom rom ( // @[Top.scala 11:21]
    .clock(rom_clock),
    .io_addr(rom_io_addr),
    .io_inst(rom_io_inst)
  );
  Ram ram ( // @[Top.scala 12:21]
    .clock(ram_clock),
    .io_addr(ram_io_addr),
    .io_rdata(ram_io_rdata),
    .io_wen(ram_io_wen),
    .io_wdata(ram_io_wdata),
    .io_rwtype(ram_io_rwtype)
  );
  Seg seg ( // @[Top.scala 13:21]
    .io_data(seg_io_data),
    .io_led_0(seg_io_led_0),
    .io_led_1(seg_io_led_1),
    .io_led_2(seg_io_led_2),
    .io_led_3(seg_io_led_3),
    .io_led_4(seg_io_led_4),
    .io_led_5(seg_io_led_5),
    .io_led_6(seg_io_led_6),
    .io_led_7(seg_io_led_7)
  );
  assign io_led_0 = seg_io_led_0; // @[Top.scala 18:12]
  assign io_led_1 = seg_io_led_1; // @[Top.scala 18:12]
  assign io_led_2 = seg_io_led_2; // @[Top.scala 18:12]
  assign io_led_3 = seg_io_led_3; // @[Top.scala 18:12]
  assign io_led_4 = seg_io_led_4; // @[Top.scala 18:12]
  assign io_led_5 = seg_io_led_5; // @[Top.scala 18:12]
  assign io_led_6 = seg_io_led_6; // @[Top.scala 18:12]
  assign io_led_7 = seg_io_led_7; // @[Top.scala 18:12]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_inst = rom_io_inst; // @[Top.scala 15:18]
  assign core_io_dmem_rdata = ram_io_rdata; // @[Top.scala 16:18]
  assign rom_clock = clock;
  assign rom_io_addr = core_io_imem_addr; // @[Top.scala 15:18]
  assign ram_clock = clock;
  assign ram_io_addr = core_io_dmem_addr; // @[Top.scala 16:18]
  assign ram_io_wen = core_io_dmem_wen; // @[Top.scala 16:18]
  assign ram_io_wdata = core_io_dmem_wdata; // @[Top.scala 16:18]
  assign ram_io_rwtype = core_io_dmem_rwtype; // @[Top.scala 16:18]
  assign seg_io_data = core_io_data; // @[Top.scala 17:18]
endmodule
